
//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/mgc_in_wire_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_wire_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule


//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.3d/815731 Production Release
//  HLS Date:       Wed Apr 24 14:54:19 PDT 2019
// 
//  Generated by:   695r48@ecegrid-thin4.ecn.purdue.edu
//  Generated date: Sat Nov 13 22:48:10 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, coeffs_rsc_z, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz, out1_rsc_dat,
      out1_rsc_triosy_lz
);
  input clk;
  input rst;
  input [511:0] coeffs_rsc_z;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;


  // Interconnect Declarations
  wire [511:0] coeffs_rsci_d;
  wire [15:0] in1_rsci_idat;
  reg [15:0] out1_rsci_idat;
  reg out1_rsc_triosy_obj_ld;
  reg main_stage_0_3;
  reg reg_in1_rsc_triosy_obj_ld_cse;
  reg [15:0] regs_1_sva;
  reg [15:0] regs_0_sva;
  reg [15:0] MAC_asn_62_itm;
  reg [15:0] MAC_asn_63_itm;
  reg [15:0] MAC_asn_64_itm;
  reg [15:0] MAC_asn_65_itm;
  reg [15:0] MAC_asn_66_itm;
  reg [15:0] MAC_asn_67_itm;
  reg [15:0] MAC_asn_68_itm;
  reg [15:0] MAC_asn_69_itm;
  reg [15:0] MAC_asn_70_itm;
  reg [15:0] MAC_asn_71_itm;
  reg [15:0] MAC_asn_72_itm;
  reg [15:0] MAC_asn_73_itm;
  reg [15:0] MAC_asn_74_itm;
  reg [15:0] MAC_asn_75_itm;
  reg [15:0] MAC_asn_76_itm;
  reg [15:0] MAC_asn_77_itm;
  reg [15:0] MAC_asn_78_itm;
  reg [15:0] MAC_asn_79_itm;
  reg [15:0] MAC_asn_80_itm;
  reg [15:0] MAC_asn_81_itm;
  reg [15:0] MAC_asn_82_itm;
  reg [15:0] MAC_asn_83_itm;
  reg [15:0] MAC_asn_84_itm;
  reg [15:0] MAC_asn_85_itm;
  reg [15:0] MAC_asn_86_itm;
  reg [15:0] MAC_asn_87_itm;
  reg [15:0] MAC_asn_88_itm;
  reg [15:0] MAC_asn_89_itm;
  reg [15:0] MAC_asn_90_itm;
  reg [29:0] MAC_acc_17_itm_1;
  wire [30:0] nl_MAC_acc_17_itm_1;
  reg [29:0] MAC_acc_16_itm_1;
  wire [30:0] nl_MAC_acc_16_itm_1;
  reg [29:0] MAC_acc_15_itm_1;
  wire [30:0] nl_MAC_acc_15_itm_1;
  reg [29:0] MAC_acc_14_itm_1;
  wire [30:0] nl_MAC_acc_14_itm_1;
  reg [29:0] MAC_acc_13_itm_1;
  wire [30:0] nl_MAC_acc_13_itm_1;
  reg [29:0] MAC_acc_12_itm_1;
  wire [30:0] nl_MAC_acc_12_itm_1;
  reg [29:0] MAC_acc_11_itm_1;
  wire [30:0] nl_MAC_acc_11_itm_1;
  reg [29:0] MAC_acc_10_itm_1;
  wire [30:0] nl_MAC_acc_10_itm_1;
  reg [29:0] MAC_acc_31_itm_1;
  wire [30:0] nl_MAC_acc_31_itm_1;
  reg [29:0] MAC_acc_9_itm_1;
  wire [30:0] nl_MAC_acc_9_itm_1;
  reg [29:0] MAC_acc_8_itm_1;
  wire [30:0] nl_MAC_acc_8_itm_1;
  reg [29:0] MAC_acc_7_itm_1;
  wire [30:0] nl_MAC_acc_7_itm_1;
  reg [29:0] MAC_acc_6_itm_1;
  wire [30:0] nl_MAC_acc_6_itm_1;
  reg [29:0] MAC_acc_5_itm_1;
  wire [30:0] nl_MAC_acc_5_itm_1;
  reg [29:0] MAC_acc_4_itm_1;
  wire [30:0] nl_MAC_acc_4_itm_1;
  reg [29:0] MAC_acc_3_itm_1;
  wire [30:0] nl_MAC_acc_3_itm_1;
  reg [29:0] MAC_acc_18_itm_1;
  wire [30:0] nl_MAC_acc_18_itm_1;
  reg [29:0] MAC_acc_itm_1;
  wire [30:0] nl_MAC_acc_itm_1;

  wire[29:0] MAC_32_acc_1_nl;
  wire[30:0] nl_MAC_32_acc_1_nl;
  wire[29:0] MAC_acc_29_nl;
  wire[30:0] nl_MAC_acc_29_nl;
  wire[29:0] MAC_acc_25_nl;
  wire[30:0] nl_MAC_acc_25_nl;
  wire[29:0] MAC_acc_24_nl;
  wire[30:0] nl_MAC_acc_24_nl;
  wire[29:0] MAC_acc_28_nl;
  wire[30:0] nl_MAC_acc_28_nl;
  wire[29:0] MAC_acc_23_nl;
  wire[30:0] nl_MAC_acc_23_nl;
  wire[29:0] MAC_acc_22_nl;
  wire[30:0] nl_MAC_acc_22_nl;
  wire[29:0] MAC_acc_27_nl;
  wire[30:0] nl_MAC_acc_27_nl;
  wire[29:0] MAC_acc_21_nl;
  wire[30:0] nl_MAC_acc_21_nl;
  wire[29:0] MAC_acc_20_nl;
  wire[30:0] nl_MAC_acc_20_nl;
  wire[29:0] MAC_acc_30_nl;
  wire[30:0] nl_MAC_acc_30_nl;
  wire[29:0] MAC_acc_19_nl;
  wire[30:0] nl_MAC_acc_19_nl;
  wire[29:0] MAC_acc_26_nl;
  wire[30:0] nl_MAC_acc_26_nl;
  wire[29:0] MAC_17_mul_nl;
  wire signed [31:0] nl_MAC_17_mul_nl;
  wire[29:0] MAC_18_mul_nl;
  wire signed [31:0] nl_MAC_18_mul_nl;
  wire[29:0] MAC_19_mul_nl;
  wire signed [31:0] nl_MAC_19_mul_nl;
  wire[29:0] MAC_20_mul_nl;
  wire signed [31:0] nl_MAC_20_mul_nl;
  wire[29:0] MAC_21_mul_nl;
  wire signed [31:0] nl_MAC_21_mul_nl;
  wire[29:0] MAC_22_mul_nl;
  wire signed [31:0] nl_MAC_22_mul_nl;
  wire[29:0] MAC_23_mul_nl;
  wire signed [31:0] nl_MAC_23_mul_nl;
  wire[29:0] MAC_24_mul_nl;
  wire signed [31:0] nl_MAC_24_mul_nl;
  wire[29:0] MAC_25_mul_nl;
  wire signed [31:0] nl_MAC_25_mul_nl;
  wire[29:0] MAC_26_mul_nl;
  wire signed [31:0] nl_MAC_26_mul_nl;
  wire[29:0] MAC_27_mul_nl;
  wire signed [31:0] nl_MAC_27_mul_nl;
  wire[29:0] MAC_28_mul_nl;
  wire signed [31:0] nl_MAC_28_mul_nl;
  wire[29:0] MAC_29_mul_nl;
  wire signed [31:0] nl_MAC_29_mul_nl;
  wire[29:0] MAC_30_mul_nl;
  wire signed [31:0] nl_MAC_30_mul_nl;
  wire[29:0] MAC_31_mul_nl;
  wire signed [31:0] nl_MAC_31_mul_nl;
  wire[29:0] MAC_32_mul_nl;
  wire signed [31:0] nl_MAC_32_mul_nl;
  wire[29:0] MAC_1_mul_nl;
  wire signed [31:0] nl_MAC_1_mul_nl;
  wire[29:0] MAC_2_mul_nl;
  wire signed [31:0] nl_MAC_2_mul_nl;
  wire[29:0] MAC_3_mul_nl;
  wire signed [31:0] nl_MAC_3_mul_nl;
  wire[29:0] MAC_4_mul_nl;
  wire signed [31:0] nl_MAC_4_mul_nl;
  wire[29:0] MAC_5_mul_nl;
  wire signed [31:0] nl_MAC_5_mul_nl;
  wire[29:0] MAC_6_mul_nl;
  wire signed [31:0] nl_MAC_6_mul_nl;
  wire[29:0] MAC_7_mul_nl;
  wire signed [31:0] nl_MAC_7_mul_nl;
  wire[29:0] MAC_8_mul_nl;
  wire signed [31:0] nl_MAC_8_mul_nl;
  wire[29:0] MAC_9_mul_nl;
  wire signed [31:0] nl_MAC_9_mul_nl;
  wire[29:0] MAC_10_mul_nl;
  wire signed [31:0] nl_MAC_10_mul_nl;
  wire[29:0] MAC_11_mul_nl;
  wire signed [31:0] nl_MAC_11_mul_nl;
  wire[29:0] MAC_12_mul_nl;
  wire signed [31:0] nl_MAC_12_mul_nl;
  wire[29:0] MAC_13_mul_nl;
  wire signed [31:0] nl_MAC_13_mul_nl;
  wire[29:0] MAC_14_mul_nl;
  wire signed [31:0] nl_MAC_14_mul_nl;
  wire[29:0] MAC_15_mul_nl;
  wire signed [31:0] nl_MAC_15_mul_nl;
  wire[29:0] MAC_16_mul_nl;
  wire signed [31:0] nl_MAC_16_mul_nl;

  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_v2 #(.rscid(32'sd1),
  .width(32'sd512)) coeffs_rsci (
      .d(coeffs_rsci_d),
      .z(coeffs_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd16)) in1_rsci (
      .dat(in1_rsc_dat),
      .idat(in1_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd16)) out1_rsci (
      .idat(out1_rsci_idat),
      .dat(out1_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) coeffs_rsc_triosy_obj (
      .ld(reg_in1_rsc_triosy_obj_ld_cse),
      .lz(coeffs_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) in1_rsc_triosy_obj (
      .ld(reg_in1_rsc_triosy_obj_ld_cse),
      .lz(in1_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) out1_rsc_triosy_obj (
      .ld(out1_rsc_triosy_obj_ld),
      .lz(out1_rsc_triosy_lz)
    );
  always @(posedge clk) begin
    if ( rst ) begin
      out1_rsc_triosy_obj_ld <= 1'b0;
      MAC_acc_31_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_itm_1 <= 30'b000000000000000000000000000000;
      reg_in1_rsc_triosy_obj_ld_cse <= 1'b0;
      main_stage_0_3 <= 1'b0;
      MAC_acc_9_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_8_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_7_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_6_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_5_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_4_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_3_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_18_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_17_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_16_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_15_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_14_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_13_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_12_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_11_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_10_itm_1 <= 30'b000000000000000000000000000000;
      MAC_asn_89_itm <= 16'b0000000000000000;
      MAC_asn_90_itm <= 16'b0000000000000000;
      MAC_asn_87_itm <= 16'b0000000000000000;
      MAC_asn_88_itm <= 16'b0000000000000000;
      MAC_asn_85_itm <= 16'b0000000000000000;
      MAC_asn_86_itm <= 16'b0000000000000000;
      MAC_asn_83_itm <= 16'b0000000000000000;
      MAC_asn_84_itm <= 16'b0000000000000000;
      MAC_asn_81_itm <= 16'b0000000000000000;
      MAC_asn_82_itm <= 16'b0000000000000000;
      MAC_asn_79_itm <= 16'b0000000000000000;
      MAC_asn_80_itm <= 16'b0000000000000000;
      MAC_asn_77_itm <= 16'b0000000000000000;
      MAC_asn_78_itm <= 16'b0000000000000000;
      MAC_asn_75_itm <= 16'b0000000000000000;
      MAC_asn_76_itm <= 16'b0000000000000000;
      MAC_asn_73_itm <= 16'b0000000000000000;
      MAC_asn_74_itm <= 16'b0000000000000000;
      MAC_asn_71_itm <= 16'b0000000000000000;
      MAC_asn_72_itm <= 16'b0000000000000000;
      MAC_asn_69_itm <= 16'b0000000000000000;
      MAC_asn_70_itm <= 16'b0000000000000000;
      MAC_asn_67_itm <= 16'b0000000000000000;
      MAC_asn_68_itm <= 16'b0000000000000000;
      MAC_asn_65_itm <= 16'b0000000000000000;
      MAC_asn_66_itm <= 16'b0000000000000000;
      MAC_asn_63_itm <= 16'b0000000000000000;
      MAC_asn_64_itm <= 16'b0000000000000000;
      regs_1_sva <= 16'b0000000000000000;
      MAC_asn_62_itm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else begin
      out1_rsc_triosy_obj_ld <= main_stage_0_3;
      MAC_acc_31_itm_1 <= nl_MAC_acc_31_itm_1[29:0];
      MAC_acc_itm_1 <= nl_MAC_acc_itm_1[29:0];
      reg_in1_rsc_triosy_obj_ld_cse <= 1'b1;
      main_stage_0_3 <= reg_in1_rsc_triosy_obj_ld_cse;
      MAC_acc_9_itm_1 <= nl_MAC_acc_9_itm_1[29:0];
      MAC_acc_8_itm_1 <= nl_MAC_acc_8_itm_1[29:0];
      MAC_acc_7_itm_1 <= nl_MAC_acc_7_itm_1[29:0];
      MAC_acc_6_itm_1 <= nl_MAC_acc_6_itm_1[29:0];
      MAC_acc_5_itm_1 <= nl_MAC_acc_5_itm_1[29:0];
      MAC_acc_4_itm_1 <= nl_MAC_acc_4_itm_1[29:0];
      MAC_acc_3_itm_1 <= nl_MAC_acc_3_itm_1[29:0];
      MAC_acc_18_itm_1 <= nl_MAC_acc_18_itm_1[29:0];
      MAC_acc_17_itm_1 <= nl_MAC_acc_17_itm_1[29:0];
      MAC_acc_16_itm_1 <= nl_MAC_acc_16_itm_1[29:0];
      MAC_acc_15_itm_1 <= nl_MAC_acc_15_itm_1[29:0];
      MAC_acc_14_itm_1 <= nl_MAC_acc_14_itm_1[29:0];
      MAC_acc_13_itm_1 <= nl_MAC_acc_13_itm_1[29:0];
      MAC_acc_12_itm_1 <= nl_MAC_acc_12_itm_1[29:0];
      MAC_acc_11_itm_1 <= nl_MAC_acc_11_itm_1[29:0];
      MAC_acc_10_itm_1 <= nl_MAC_acc_10_itm_1[29:0];
      MAC_asn_89_itm <= MAC_asn_88_itm;
      MAC_asn_90_itm <= MAC_asn_89_itm;
      MAC_asn_87_itm <= MAC_asn_86_itm;
      MAC_asn_88_itm <= MAC_asn_87_itm;
      MAC_asn_85_itm <= MAC_asn_84_itm;
      MAC_asn_86_itm <= MAC_asn_85_itm;
      MAC_asn_83_itm <= MAC_asn_82_itm;
      MAC_asn_84_itm <= MAC_asn_83_itm;
      MAC_asn_81_itm <= MAC_asn_80_itm;
      MAC_asn_82_itm <= MAC_asn_81_itm;
      MAC_asn_79_itm <= MAC_asn_78_itm;
      MAC_asn_80_itm <= MAC_asn_79_itm;
      MAC_asn_77_itm <= MAC_asn_76_itm;
      MAC_asn_78_itm <= MAC_asn_77_itm;
      MAC_asn_75_itm <= MAC_asn_74_itm;
      MAC_asn_76_itm <= MAC_asn_75_itm;
      MAC_asn_73_itm <= MAC_asn_72_itm;
      MAC_asn_74_itm <= MAC_asn_73_itm;
      MAC_asn_71_itm <= MAC_asn_70_itm;
      MAC_asn_72_itm <= MAC_asn_71_itm;
      MAC_asn_69_itm <= MAC_asn_68_itm;
      MAC_asn_70_itm <= MAC_asn_69_itm;
      MAC_asn_67_itm <= MAC_asn_66_itm;
      MAC_asn_68_itm <= MAC_asn_67_itm;
      MAC_asn_65_itm <= MAC_asn_64_itm;
      MAC_asn_66_itm <= MAC_asn_65_itm;
      MAC_asn_63_itm <= MAC_asn_62_itm;
      MAC_asn_64_itm <= MAC_asn_63_itm;
      regs_1_sva <= regs_0_sva;
      MAC_asn_62_itm <= regs_1_sva;
      regs_0_sva <= in1_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out1_rsci_idat <= 16'b0000000000000000;
    end
    else if ( main_stage_0_3 ) begin
      out1_rsci_idat <= readslicef_30_16_14((MAC_32_acc_1_nl));
    end
  end
  assign nl_MAC_acc_25_nl = MAC_acc_17_itm_1 + MAC_acc_16_itm_1;
  assign MAC_acc_25_nl = nl_MAC_acc_25_nl[29:0];
  assign nl_MAC_acc_24_nl = MAC_acc_15_itm_1 + MAC_acc_14_itm_1;
  assign MAC_acc_24_nl = nl_MAC_acc_24_nl[29:0];
  assign nl_MAC_acc_29_nl = (MAC_acc_25_nl) + (MAC_acc_24_nl);
  assign MAC_acc_29_nl = nl_MAC_acc_29_nl[29:0];
  assign nl_MAC_acc_23_nl = MAC_acc_13_itm_1 + MAC_acc_12_itm_1;
  assign MAC_acc_23_nl = nl_MAC_acc_23_nl[29:0];
  assign nl_MAC_acc_22_nl = MAC_acc_11_itm_1 + MAC_acc_10_itm_1;
  assign MAC_acc_22_nl = nl_MAC_acc_22_nl[29:0];
  assign nl_MAC_acc_28_nl = (MAC_acc_23_nl) + (MAC_acc_22_nl);
  assign MAC_acc_28_nl = nl_MAC_acc_28_nl[29:0];
  assign nl_MAC_acc_31_itm_1  = (MAC_acc_29_nl) + (MAC_acc_28_nl);
  assign nl_MAC_acc_21_nl = MAC_acc_9_itm_1 + MAC_acc_8_itm_1;
  assign MAC_acc_21_nl = nl_MAC_acc_21_nl[29:0];
  assign nl_MAC_acc_20_nl = MAC_acc_7_itm_1 + MAC_acc_6_itm_1;
  assign MAC_acc_20_nl = nl_MAC_acc_20_nl[29:0];
  assign nl_MAC_acc_27_nl = (MAC_acc_21_nl) + (MAC_acc_20_nl);
  assign MAC_acc_27_nl = nl_MAC_acc_27_nl[29:0];
  assign nl_MAC_acc_19_nl = MAC_acc_5_itm_1 + MAC_acc_4_itm_1;
  assign MAC_acc_19_nl = nl_MAC_acc_19_nl[29:0];
  assign nl_MAC_acc_26_nl = MAC_acc_3_itm_1 + MAC_acc_18_itm_1;
  assign MAC_acc_26_nl = nl_MAC_acc_26_nl[29:0];
  assign nl_MAC_acc_30_nl = (MAC_acc_19_nl) + (MAC_acc_26_nl);
  assign MAC_acc_30_nl = nl_MAC_acc_30_nl[29:0];
  assign nl_MAC_acc_itm_1  = (MAC_acc_27_nl) + (MAC_acc_30_nl);
  assign nl_MAC_17_mul_nl = $signed(MAC_asn_75_itm) * $signed((coeffs_rsci_d[271:256]));
  assign MAC_17_mul_nl = nl_MAC_17_mul_nl[29:0];
  assign nl_MAC_18_mul_nl = $signed(MAC_asn_76_itm) * $signed((coeffs_rsci_d[287:272]));
  assign MAC_18_mul_nl = nl_MAC_18_mul_nl[29:0];
  assign nl_MAC_acc_9_itm_1  = (MAC_17_mul_nl) + (MAC_18_mul_nl);
  assign nl_MAC_19_mul_nl = $signed(MAC_asn_77_itm) * $signed((coeffs_rsci_d[303:288]));
  assign MAC_19_mul_nl = nl_MAC_19_mul_nl[29:0];
  assign nl_MAC_20_mul_nl = $signed(MAC_asn_78_itm) * $signed((coeffs_rsci_d[319:304]));
  assign MAC_20_mul_nl = nl_MAC_20_mul_nl[29:0];
  assign nl_MAC_acc_8_itm_1  = (MAC_19_mul_nl) + (MAC_20_mul_nl);
  assign nl_MAC_21_mul_nl = $signed(MAC_asn_79_itm) * $signed((coeffs_rsci_d[335:320]));
  assign MAC_21_mul_nl = nl_MAC_21_mul_nl[29:0];
  assign nl_MAC_22_mul_nl = $signed(MAC_asn_80_itm) * $signed((coeffs_rsci_d[351:336]));
  assign MAC_22_mul_nl = nl_MAC_22_mul_nl[29:0];
  assign nl_MAC_acc_7_itm_1  = (MAC_21_mul_nl) + (MAC_22_mul_nl);
  assign nl_MAC_23_mul_nl = $signed(MAC_asn_81_itm) * $signed((coeffs_rsci_d[367:352]));
  assign MAC_23_mul_nl = nl_MAC_23_mul_nl[29:0];
  assign nl_MAC_24_mul_nl = $signed(MAC_asn_82_itm) * $signed((coeffs_rsci_d[383:368]));
  assign MAC_24_mul_nl = nl_MAC_24_mul_nl[29:0];
  assign nl_MAC_acc_6_itm_1  = (MAC_23_mul_nl) + (MAC_24_mul_nl);
  assign nl_MAC_25_mul_nl = $signed(MAC_asn_83_itm) * $signed((coeffs_rsci_d[399:384]));
  assign MAC_25_mul_nl = nl_MAC_25_mul_nl[29:0];
  assign nl_MAC_26_mul_nl = $signed(MAC_asn_84_itm) * $signed((coeffs_rsci_d[415:400]));
  assign MAC_26_mul_nl = nl_MAC_26_mul_nl[29:0];
  assign nl_MAC_acc_5_itm_1  = (MAC_25_mul_nl) + (MAC_26_mul_nl);
  assign nl_MAC_27_mul_nl = $signed(MAC_asn_85_itm) * $signed((coeffs_rsci_d[431:416]));
  assign MAC_27_mul_nl = nl_MAC_27_mul_nl[29:0];
  assign nl_MAC_28_mul_nl = $signed(MAC_asn_86_itm) * $signed((coeffs_rsci_d[447:432]));
  assign MAC_28_mul_nl = nl_MAC_28_mul_nl[29:0];
  assign nl_MAC_acc_4_itm_1  = (MAC_27_mul_nl) + (MAC_28_mul_nl);
  assign nl_MAC_29_mul_nl = $signed(MAC_asn_87_itm) * $signed((coeffs_rsci_d[463:448]));
  assign MAC_29_mul_nl = nl_MAC_29_mul_nl[29:0];
  assign nl_MAC_30_mul_nl = $signed(MAC_asn_88_itm) * $signed((coeffs_rsci_d[479:464]));
  assign MAC_30_mul_nl = nl_MAC_30_mul_nl[29:0];
  assign nl_MAC_acc_3_itm_1  = (MAC_29_mul_nl) + (MAC_30_mul_nl);
  assign nl_MAC_31_mul_nl = $signed(MAC_asn_89_itm) * $signed((coeffs_rsci_d[495:480]));
  assign MAC_31_mul_nl = nl_MAC_31_mul_nl[29:0];
  assign nl_MAC_32_mul_nl = $signed(MAC_asn_90_itm) * $signed((coeffs_rsci_d[511:496]));
  assign MAC_32_mul_nl = nl_MAC_32_mul_nl[29:0];
  assign nl_MAC_acc_18_itm_1  = (MAC_31_mul_nl) + (MAC_32_mul_nl);
  assign nl_MAC_1_mul_nl = $signed((in1_rsci_idat)) * $signed((coeffs_rsci_d[15:0]));
  assign MAC_1_mul_nl = nl_MAC_1_mul_nl[29:0];
  assign nl_MAC_2_mul_nl = $signed(regs_0_sva) * $signed((coeffs_rsci_d[31:16]));
  assign MAC_2_mul_nl = nl_MAC_2_mul_nl[29:0];
  assign nl_MAC_acc_17_itm_1  = (MAC_1_mul_nl) + (MAC_2_mul_nl);
  assign nl_MAC_3_mul_nl = $signed(regs_1_sva) * $signed((coeffs_rsci_d[47:32]));
  assign MAC_3_mul_nl = nl_MAC_3_mul_nl[29:0];
  assign nl_MAC_4_mul_nl = $signed(MAC_asn_62_itm) * $signed((coeffs_rsci_d[63:48]));
  assign MAC_4_mul_nl = nl_MAC_4_mul_nl[29:0];
  assign nl_MAC_acc_16_itm_1  = (MAC_3_mul_nl) + (MAC_4_mul_nl);
  assign nl_MAC_5_mul_nl = $signed(MAC_asn_63_itm) * $signed((coeffs_rsci_d[79:64]));
  assign MAC_5_mul_nl = nl_MAC_5_mul_nl[29:0];
  assign nl_MAC_6_mul_nl = $signed(MAC_asn_64_itm) * $signed((coeffs_rsci_d[95:80]));
  assign MAC_6_mul_nl = nl_MAC_6_mul_nl[29:0];
  assign nl_MAC_acc_15_itm_1  = (MAC_5_mul_nl) + (MAC_6_mul_nl);
  assign nl_MAC_7_mul_nl = $signed(MAC_asn_65_itm) * $signed((coeffs_rsci_d[111:96]));
  assign MAC_7_mul_nl = nl_MAC_7_mul_nl[29:0];
  assign nl_MAC_8_mul_nl = $signed(MAC_asn_66_itm) * $signed((coeffs_rsci_d[127:112]));
  assign MAC_8_mul_nl = nl_MAC_8_mul_nl[29:0];
  assign nl_MAC_acc_14_itm_1  = (MAC_7_mul_nl) + (MAC_8_mul_nl);
  assign nl_MAC_9_mul_nl = $signed(MAC_asn_67_itm) * $signed((coeffs_rsci_d[143:128]));
  assign MAC_9_mul_nl = nl_MAC_9_mul_nl[29:0];
  assign nl_MAC_10_mul_nl = $signed(MAC_asn_68_itm) * $signed((coeffs_rsci_d[159:144]));
  assign MAC_10_mul_nl = nl_MAC_10_mul_nl[29:0];
  assign nl_MAC_acc_13_itm_1  = (MAC_9_mul_nl) + (MAC_10_mul_nl);
  assign nl_MAC_11_mul_nl = $signed(MAC_asn_69_itm) * $signed((coeffs_rsci_d[175:160]));
  assign MAC_11_mul_nl = nl_MAC_11_mul_nl[29:0];
  assign nl_MAC_12_mul_nl = $signed(MAC_asn_70_itm) * $signed((coeffs_rsci_d[191:176]));
  assign MAC_12_mul_nl = nl_MAC_12_mul_nl[29:0];
  assign nl_MAC_acc_12_itm_1  = (MAC_11_mul_nl) + (MAC_12_mul_nl);
  assign nl_MAC_13_mul_nl = $signed(MAC_asn_71_itm) * $signed((coeffs_rsci_d[207:192]));
  assign MAC_13_mul_nl = nl_MAC_13_mul_nl[29:0];
  assign nl_MAC_14_mul_nl = $signed(MAC_asn_72_itm) * $signed((coeffs_rsci_d[223:208]));
  assign MAC_14_mul_nl = nl_MAC_14_mul_nl[29:0];
  assign nl_MAC_acc_11_itm_1  = (MAC_13_mul_nl) + (MAC_14_mul_nl);
  assign nl_MAC_15_mul_nl = $signed(MAC_asn_73_itm) * $signed((coeffs_rsci_d[239:224]));
  assign MAC_15_mul_nl = nl_MAC_15_mul_nl[29:0];
  assign nl_MAC_16_mul_nl = $signed(MAC_asn_74_itm) * $signed((coeffs_rsci_d[255:240]));
  assign MAC_16_mul_nl = nl_MAC_16_mul_nl[29:0];
  assign nl_MAC_acc_10_itm_1  = (MAC_15_mul_nl) + (MAC_16_mul_nl);
  assign nl_MAC_32_acc_1_nl = MAC_acc_31_itm_1 + MAC_acc_itm_1;
  assign MAC_32_acc_1_nl = nl_MAC_32_acc_1_nl[29:0];

  function automatic [15:0] readslicef_30_16_14;
    input [29:0] vector;
    reg [29:0] tmp;
  begin
    tmp = vector >> 14;
    readslicef_30_16_14 = tmp[15:0];
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, coeffs_rsc_z, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz, out1_rsc_dat,
      out1_rsc_triosy_lz
);
  input clk;
  input rst;
  input [511:0] coeffs_rsc_z;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .coeffs_rsc_z(coeffs_rsc_z),
      .coeffs_rsc_triosy_lz(coeffs_rsc_triosy_lz),
      .in1_rsc_dat(in1_rsc_dat),
      .in1_rsc_triosy_lz(in1_rsc_triosy_lz),
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_triosy_lz(out1_rsc_triosy_lz)
    );
endmodule



