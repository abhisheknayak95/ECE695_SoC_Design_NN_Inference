
--------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_out_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_out_pkg_v1 IS

COMPONENT ccs_out_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    dat    : OUT std_logic_vector(width-1 DOWNTO 0);
    idat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_out_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_out_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    dat   : OUT std_logic_vector(width-1 DOWNTO 0);
    idat  : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_out_v1;

ARCHITECTURE beh OF ccs_out_v1 IS
BEGIN

  dat <= idat;

END beh;


--------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.3d/815731 Production Release
--  HLS Date:       Wed Apr 24 14:54:19 PDT 2019
-- 
--  Generated by:   695r48@cparch23.ecn.purdue.edu
--  Generated date: Tue Nov  9 16:00:03 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen IS
  PORT(
    q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    rport_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen;

ARCHITECTURE v14 OF fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen IS
  -- Default Constants

BEGIN
  q_d <= q;
  radr <= (radr_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    fir_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY fir_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (34 DOWNTO 0)
  );
END fir_core_core_fsm;

ARCHITECTURE v14 OF fir_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for fir_core_core_fsm_1
  TYPE fir_core_core_fsm_1_ST IS (core_rlp_C_0, main_C_0, main_C_1, main_C_2, main_C_3,
      main_C_4, main_C_5, main_C_6, main_C_7, main_C_8, main_C_9, main_C_10, main_C_11,
      main_C_12, main_C_13, main_C_14, main_C_15, main_C_16, main_C_17, main_C_18,
      main_C_19, main_C_20, main_C_21, main_C_22, main_C_23, main_C_24, main_C_25,
      main_C_26, main_C_27, main_C_28, main_C_29, main_C_30, main_C_31, main_C_32,
      main_C_33);

  SIGNAL state_var : fir_core_core_fsm_1_ST;
  SIGNAL state_var_NS : fir_core_core_fsm_1_ST;

BEGIN
  fir_core_core_fsm_1 : PROCESS (state_var)
  BEGIN
    CASE state_var IS
      WHEN main_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000010");
        state_var_NS <= main_C_1;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000100");
        state_var_NS <= main_C_2;
      WHEN main_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000001000");
        state_var_NS <= main_C_3;
      WHEN main_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000010000");
        state_var_NS <= main_C_4;
      WHEN main_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000100000");
        state_var_NS <= main_C_5;
      WHEN main_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000001000000");
        state_var_NS <= main_C_6;
      WHEN main_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000010000000");
        state_var_NS <= main_C_7;
      WHEN main_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000100000000");
        state_var_NS <= main_C_8;
      WHEN main_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000001000000000");
        state_var_NS <= main_C_9;
      WHEN main_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000010000000000");
        state_var_NS <= main_C_10;
      WHEN main_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000100000000000");
        state_var_NS <= main_C_11;
      WHEN main_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000001000000000000");
        state_var_NS <= main_C_12;
      WHEN main_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000010000000000000");
        state_var_NS <= main_C_13;
      WHEN main_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000100000000000000");
        state_var_NS <= main_C_14;
      WHEN main_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000001000000000000000");
        state_var_NS <= main_C_15;
      WHEN main_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000010000000000000000");
        state_var_NS <= main_C_16;
      WHEN main_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000100000000000000000");
        state_var_NS <= main_C_17;
      WHEN main_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000001000000000000000000");
        state_var_NS <= main_C_18;
      WHEN main_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000010000000000000000000");
        state_var_NS <= main_C_19;
      WHEN main_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000100000000000000000000");
        state_var_NS <= main_C_20;
      WHEN main_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000001000000000000000000000");
        state_var_NS <= main_C_21;
      WHEN main_C_21 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000010000000000000000000000");
        state_var_NS <= main_C_22;
      WHEN main_C_22 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000100000000000000000000000");
        state_var_NS <= main_C_23;
      WHEN main_C_23 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000001000000000000000000000000");
        state_var_NS <= main_C_24;
      WHEN main_C_24 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000010000000000000000000000000");
        state_var_NS <= main_C_25;
      WHEN main_C_25 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000100000000000000000000000000");
        state_var_NS <= main_C_26;
      WHEN main_C_26 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001000000000000000000000000000");
        state_var_NS <= main_C_27;
      WHEN main_C_27 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010000000000000000000000000000");
        state_var_NS <= main_C_28;
      WHEN main_C_28 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100000000000000000000000000000");
        state_var_NS <= main_C_29;
      WHEN main_C_29 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000000000000000000000000000000");
        state_var_NS <= main_C_30;
      WHEN main_C_30 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000000000000000000000000000000");
        state_var_NS <= main_C_31;
      WHEN main_C_31 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000000000000000000000000000000");
        state_var_NS <= main_C_32;
      WHEN main_C_32 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000000000000000000000000000000");
        state_var_NS <= main_C_33;
      WHEN main_C_33 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000000000000000000000000000000");
        state_var_NS <= main_C_0;
      -- core_rlp_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000001");
        state_var_NS <= main_C_0;
    END CASE;
  END PROCESS fir_core_core_fsm_1;

  fir_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= core_rlp_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS fir_core_core_fsm_1_REG;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    fir_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY fir_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    coeffs_rsc_triosy_lz : OUT STD_LOGIC;
    in1_rsc_dat : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    in1_rsc_triosy_lz : OUT STD_LOGIC;
    out1_rsc_dat : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    out1_rsc_triosy_lz : OUT STD_LOGIC;
    coeffs_rsci_radr_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    coeffs_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC
  );
END fir_core;

ARCHITECTURE v14 OF fir_core IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL in1_rsci_idat : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL out1_rsci_idat : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL coeffs_rsc_triosy_obj_ld : STD_LOGIC;
  SIGNAL in1_rsc_triosy_obj_ld : STD_LOGIC;
  SIGNAL out1_rsc_triosy_obj_ld : STD_LOGIC;
  SIGNAL fsm_output : STD_LOGIC_VECTOR (34 DOWNTO 0);
  SIGNAL main_stage_0_2 : STD_LOGIC;
  SIGNAL reg_MAC_asn_89_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_88_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_87_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_86_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_85_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_84_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_83_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_82_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_81_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_80_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_79_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_78_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_77_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_76_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_75_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_74_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_73_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_72_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_71_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_70_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_69_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_68_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_67_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_66_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_65_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_64_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL reg_MAC_asn_63_cse : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL z_out : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL regs_3_sva : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL regs_2_sva : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL regs_0_sva : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL asn_ncse_sva : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_asn_62_itm : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_10_mul_itm : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_11_mul_itm : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_10_itm : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_22_itm : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_28_itm : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_asn_90_itm : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL MAC_acc_itm : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_28_itm_mx0w17 : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_31_mx0w0 : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_26_itm_mx0w1 : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_10_itm_mx0c0 : STD_LOGIC;
  SIGNAL MAC_acc_10_itm_mx0c1 : STD_LOGIC;
  SIGNAL MAC_acc_22_itm_mx0c2 : STD_LOGIC;

  SIGNAL MAC_32_acc_1_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_32_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_30_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_28_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_26_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_24_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_22_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_20_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_18_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_16_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_14_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_12_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_10_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_8_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_6_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_4_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_2_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_31_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_29_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_27_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_25_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_23_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_21_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_19_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_17_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_27_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_21_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_15_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_13_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_11_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_9_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_7_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_5_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_3_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_1_mul_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL MAC_acc_30_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL mux1h_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL coeffs_nor_nl : STD_LOGIC;
  SIGNAL MAC_mux_2_nl : STD_LOGIC_VECTOR (29 DOWNTO 0);
  SIGNAL in1_rsci_dat : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL in1_rsci_idat_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  SIGNAL out1_rsci_idat_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL out1_rsci_dat : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT fir_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (34 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL fir_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (34 DOWNTO 0);

  FUNCTION MUX1HOT_v_30_17_2(input_16 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(16 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(29 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(29 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_30_18_2(input_17 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(17 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(29 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(29 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_30_3_2(input_2 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(29 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(29 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_30_2(input_29 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(29 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_v_16_2_2(input_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(15 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_30_2_2(input_0 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(29 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  in1_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 16
      )
    PORT MAP(
      dat => in1_rsci_dat,
      idat => in1_rsci_idat_1
    );
  in1_rsci_dat <= in1_rsc_dat;
  in1_rsci_idat <= in1_rsci_idat_1;

  out1_rsci : work.ccs_out_pkg_v1.ccs_out_v1
    GENERIC MAP(
      rscid => 3,
      width => 16
      )
    PORT MAP(
      idat => out1_rsci_idat_1,
      dat => out1_rsci_dat
    );
  out1_rsci_idat_1 <= out1_rsci_idat;
  out1_rsc_dat <= out1_rsci_dat;

  coeffs_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => coeffs_rsc_triosy_obj_ld,
      lz => coeffs_rsc_triosy_lz
    );
  in1_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => in1_rsc_triosy_obj_ld,
      lz => in1_rsc_triosy_lz
    );
  out1_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => out1_rsc_triosy_obj_ld,
      lz => out1_rsc_triosy_lz
    );
  fir_core_core_fsm_inst : fir_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      fsm_output => fir_core_core_fsm_inst_fsm_output
    );
  fsm_output <= fir_core_core_fsm_inst_fsm_output;

  MAC_acc_28_itm_mx0w17 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_acc_26_itm_mx0w1)
      + UNSIGNED(MAC_acc_22_itm), 30));
  MAC_acc_31_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_11_mul_itm) + UNSIGNED(MAC_10_mul_itm),
      30));
  MAC_acc_26_itm_mx0w1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_acc_31_mx0w0)
      + UNSIGNED(MAC_acc_10_itm), 30));
  MAC_acc_10_itm_mx0c0 <= (fsm_output(28)) OR (fsm_output(24)) OR (fsm_output(20))
      OR (fsm_output(12)) OR (fsm_output(4)) OR (fsm_output(32));
  MAC_acc_10_itm_mx0c1 <= (fsm_output(14)) OR (fsm_output(6));
  MAC_acc_22_itm_mx0c2 <= (fsm_output(30)) OR (fsm_output(22));
  mux1h_nl <= MUX1HOT_v_5_30_2(STD_LOGIC_VECTOR'( "11110"), STD_LOGIC_VECTOR'( "11101"),
      STD_LOGIC_VECTOR'( "11100"), STD_LOGIC_VECTOR'( "11011"), STD_LOGIC_VECTOR'(
      "11010"), STD_LOGIC_VECTOR'( "11001"), STD_LOGIC_VECTOR'( "11000"), STD_LOGIC_VECTOR'(
      "10111"), STD_LOGIC_VECTOR'( "10110"), STD_LOGIC_VECTOR'( "10101"), STD_LOGIC_VECTOR'(
      "10100"), STD_LOGIC_VECTOR'( "10011"), STD_LOGIC_VECTOR'( "10010"), STD_LOGIC_VECTOR'(
      "10001"), STD_LOGIC_VECTOR'( "10000"), STD_LOGIC_VECTOR'( "01111"), STD_LOGIC_VECTOR'(
      "01110"), STD_LOGIC_VECTOR'( "01101"), STD_LOGIC_VECTOR'( "01100"), STD_LOGIC_VECTOR'(
      "01011"), STD_LOGIC_VECTOR'( "01010"), STD_LOGIC_VECTOR'( "01001"), STD_LOGIC_VECTOR'(
      "01000"), STD_LOGIC_VECTOR'( "00111"), STD_LOGIC_VECTOR'( "00110"), STD_LOGIC_VECTOR'(
      "00101"), STD_LOGIC_VECTOR'( "00100"), STD_LOGIC_VECTOR'( "00011"), STD_LOGIC_VECTOR'(
      "00010"), STD_LOGIC_VECTOR'( "00001"), STD_LOGIC_VECTOR'( (fsm_output(2)) &
      (fsm_output(3)) & (fsm_output(4)) & (fsm_output(5)) & (fsm_output(6)) & (fsm_output(7))
      & (fsm_output(8)) & (fsm_output(9)) & (fsm_output(10)) & (fsm_output(11)) &
      (fsm_output(12)) & (fsm_output(13)) & (fsm_output(14)) & (fsm_output(15)) &
      (fsm_output(16)) & (fsm_output(17)) & (fsm_output(18)) & (fsm_output(19)) &
      (fsm_output(20)) & (fsm_output(21)) & (fsm_output(22)) & (fsm_output(23)) &
      (fsm_output(24)) & (fsm_output(25)) & (fsm_output(26)) & (fsm_output(27)) &
      (fsm_output(28)) & (fsm_output(29)) & (fsm_output(30)) & (fsm_output(31))));
  coeffs_nor_nl <= NOT((fsm_output(0)) OR (fsm_output(33)) OR (fsm_output(34)) OR
      (fsm_output(32)));
  and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), mux1h_nl, coeffs_nor_nl);
  coeffs_rsci_radr_d <= MUX_v_5_2_2(and_nl, STD_LOGIC_VECTOR'("11111"), (fsm_output(1)));
  coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d <= NOT((fsm_output(0)) OR (fsm_output(33))
      OR (fsm_output(34)));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        out1_rsc_triosy_obj_ld <= '0';
        in1_rsc_triosy_obj_ld <= '0';
        coeffs_rsc_triosy_obj_ld <= '0';
        main_stage_0_2 <= '0';
        MAC_11_mul_itm <= STD_LOGIC_VECTOR'( "000000000000000000000000000000");
      ELSE
        out1_rsc_triosy_obj_ld <= main_stage_0_2;
        in1_rsc_triosy_obj_ld <= fsm_output(1);
        coeffs_rsc_triosy_obj_ld <= fsm_output(32);
        main_stage_0_2 <= fsm_output(34);
        MAC_11_mul_itm <= MUX1HOT_v_30_18_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_31_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_29_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_27_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_25_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_23_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_21_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_19_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_17_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_acc_27_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_15_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_13_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_11_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_9_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_7_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_5_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_3_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_1_mul_nl),
            30)), MAC_acc_28_itm_mx0w17, STD_LOGIC_VECTOR'( (fsm_output(3)) & (fsm_output(5))
            & (fsm_output(7)) & (fsm_output(9)) & (fsm_output(11)) & (fsm_output(13))
            & (fsm_output(15)) & (fsm_output(17)) & (fsm_output(18)) & (fsm_output(19))
            & (fsm_output(21)) & (fsm_output(23)) & (fsm_output(25)) & (fsm_output(27))
            & (fsm_output(29)) & (fsm_output(31)) & (fsm_output(33)) & (fsm_output(34))));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        out1_rsci_idat <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( main_stage_0_2 = '1' ) THEN
        out1_rsci_idat <= MAC_32_acc_1_nl(29 DOWNTO 14);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        regs_0_sva <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(33)) = '1' ) THEN
        regs_0_sva <= asn_ncse_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        regs_2_sva <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        regs_2_sva <= MAC_asn_62_itm;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MAC_asn_62_itm <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( ((fsm_output(34)) OR (fsm_output(32))) = '1' ) THEN
        MAC_asn_62_itm <= MUX_v_16_2_2(regs_0_sva, regs_2_sva, fsm_output(34));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_63_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_63_cse <= regs_3_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_64_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_64_cse <= reg_MAC_asn_63_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_65_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_65_cse <= reg_MAC_asn_64_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_66_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_66_cse <= reg_MAC_asn_65_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_67_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_67_cse <= reg_MAC_asn_66_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_68_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_68_cse <= reg_MAC_asn_67_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_69_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_69_cse <= reg_MAC_asn_68_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_70_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_70_cse <= reg_MAC_asn_69_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_71_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_71_cse <= reg_MAC_asn_70_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_72_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_72_cse <= reg_MAC_asn_71_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_73_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_73_cse <= reg_MAC_asn_72_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_74_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_74_cse <= reg_MAC_asn_73_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_75_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_75_cse <= reg_MAC_asn_74_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_76_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_76_cse <= reg_MAC_asn_75_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_77_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_77_cse <= reg_MAC_asn_76_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_78_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_78_cse <= reg_MAC_asn_77_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_79_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_79_cse <= reg_MAC_asn_78_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_80_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_80_cse <= reg_MAC_asn_79_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_81_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_81_cse <= reg_MAC_asn_80_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_82_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_82_cse <= reg_MAC_asn_81_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_83_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_83_cse <= reg_MAC_asn_82_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_84_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_84_cse <= reg_MAC_asn_83_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_85_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_85_cse <= reg_MAC_asn_84_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_86_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_86_cse <= reg_MAC_asn_85_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_87_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_87_cse <= reg_MAC_asn_86_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_88_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_88_cse <= reg_MAC_asn_87_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_MAC_asn_89_cse <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        reg_MAC_asn_89_cse <= reg_MAC_asn_88_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MAC_asn_90_itm <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        MAC_asn_90_itm <= reg_MAC_asn_89_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        regs_3_sva <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(34)) = '1' ) THEN
        regs_3_sva <= regs_2_sva;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MAC_10_mul_itm <= STD_LOGIC_VECTOR'( "000000000000000000000000000000");
      ELSIF ( ((fsm_output(34)) OR (fsm_output(30)) OR (fsm_output(26)) OR (fsm_output(18))
          OR (fsm_output(2)) OR (fsm_output(14)) OR (fsm_output(28)) OR (fsm_output(10))
          OR (fsm_output(8)) OR (fsm_output(22)) OR (fsm_output(16)) OR (fsm_output(4))
          OR (fsm_output(6)) OR (fsm_output(12)) OR (fsm_output(20)) OR (fsm_output(24))
          OR (fsm_output(32))) = '1' ) THEN
        MAC_10_mul_itm <= MUX1HOT_v_30_17_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_32_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_30_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_28_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_26_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_24_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_22_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_20_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_18_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_16_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_14_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_12_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_10_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_8_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_6_mul_nl), 30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_4_mul_nl),
            30)), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_2_mul_nl), 30)), MAC_acc_28_itm,
            STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6))
            & (fsm_output(8)) & (fsm_output(10)) & (fsm_output(12)) & (fsm_output(14))
            & (fsm_output(16)) & (fsm_output(18)) & (fsm_output(20)) & (fsm_output(22))
            & (fsm_output(24)) & (fsm_output(26)) & (fsm_output(28)) & (fsm_output(30))
            & (fsm_output(32)) & (fsm_output(34))));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MAC_acc_10_itm <= STD_LOGIC_VECTOR'( "000000000000000000000000000000");
      ELSIF ( (MAC_acc_10_itm_mx0c0 OR MAC_acc_10_itm_mx0c1 OR (fsm_output(34)))
          = '1' ) THEN
        MAC_acc_10_itm <= MUX1HOT_v_30_3_2(MAC_acc_31_mx0w0, MAC_acc_26_itm_mx0w1,
            MAC_acc_itm, STD_LOGIC_VECTOR'( MAC_acc_10_itm_mx0c0 & MAC_acc_10_itm_mx0c1
            & (fsm_output(34))));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        asn_ncse_sva <= STD_LOGIC_VECTOR'( "0000000000000000");
      ELSIF ( (fsm_output(1)) = '1' ) THEN
        asn_ncse_sva <= in1_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MAC_acc_22_itm <= STD_LOGIC_VECTOR'( "000000000000000000000000000000");
      ELSIF ( ((fsm_output(10)) OR (fsm_output(8)) OR MAC_acc_22_itm_mx0c2) = '1'
          ) THEN
        MAC_acc_22_itm <= MUX1HOT_v_30_3_2(MAC_acc_31_mx0w0, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_acc_30_nl),
            30)), MAC_acc_26_itm_mx0w1, STD_LOGIC_VECTOR'( (fsm_output(8)) & (fsm_output(10))
            & MAC_acc_22_itm_mx0c2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MAC_acc_28_itm <= STD_LOGIC_VECTOR'( "000000000000000000000000000000");
      ELSIF ( ((fsm_output(26)) OR (fsm_output(16))) = '1' ) THEN
        MAC_acc_28_itm <= MUX_v_30_2_2(MAC_acc_31_mx0w0, MAC_acc_28_itm_mx0w17, fsm_output(26));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        MAC_acc_itm <= STD_LOGIC_VECTOR'( "000000000000000000000000000000");
      ELSIF ( (fsm_output(19)) = '1' ) THEN
        MAC_acc_itm <= z_out;
      END IF;
    END IF;
  END PROCESS;
  MAC_31_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_89_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_29_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_87_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_27_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_85_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_25_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_83_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_23_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_81_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_21_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_79_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_19_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_77_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_17_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_75_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_acc_21_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_acc_31_mx0w0) + UNSIGNED(MAC_acc_28_itm),
      30));
  MAC_acc_27_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(MAC_acc_21_nl),
      30) + UNSIGNED(MAC_acc_10_itm), 30));
  MAC_15_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_73_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_13_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_71_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_11_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_69_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_9_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_67_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_7_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_65_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_5_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_63_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_3_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(regs_2_sva) * SIGNED(coeffs_rsci_q_d)),
      30));
  MAC_1_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(asn_ncse_sva) *
      SIGNED(coeffs_rsci_q_d)), 30));
  MAC_32_acc_1_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(MAC_acc_31_mx0w0) + SIGNED(MAC_acc_10_itm),
      30));
  MAC_32_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(MAC_asn_90_itm)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_30_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_88_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_28_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_86_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_26_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_84_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_24_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_82_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_22_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_80_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_20_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_78_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_18_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_76_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_16_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_74_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_14_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_72_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_12_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_70_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_10_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_68_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_8_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_66_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_6_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(reg_MAC_asn_64_cse)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_4_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(MAC_asn_62_itm)
      * SIGNED(coeffs_rsci_q_d)), 30));
  MAC_2_mul_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(SIGNED'( SIGNED(regs_0_sva) * SIGNED(coeffs_rsci_q_d)),
      30));
  MAC_acc_30_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(z_out) + UNSIGNED(MAC_acc_10_itm),
      30));
  MAC_mux_2_nl <= MUX_v_30_2_2(MAC_acc_31_mx0w0, MAC_11_mul_itm, fsm_output(19));
  z_out <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(MAC_mux_2_nl) + UNSIGNED(MAC_acc_22_itm),
      30));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    fir
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.ccs_in_pkg_v1.ALL;
USE work.ccs_out_pkg_v1.ALL;
USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY fir IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    coeffs_rsc_radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    coeffs_rsc_q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    coeffs_rsc_triosy_lz : OUT STD_LOGIC;
    in1_rsc_dat : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
    in1_rsc_triosy_lz : OUT STD_LOGIC;
    out1_rsc_dat : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
    out1_rsc_triosy_lz : OUT STD_LOGIC
  );
END fir;

ARCHITECTURE v14 OF fir IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL coeffs_rsci_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL coeffs_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;

  COMPONENT fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen
    PORT(
      q : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      radr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      q_d : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      rport_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL coeffs_rsci_q : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL coeffs_rsci_radr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL coeffs_rsci_radr_d_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL coeffs_rsci_q_d_1 : STD_LOGIC_VECTOR (15 DOWNTO 0);

  COMPONENT fir_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      coeffs_rsc_triosy_lz : OUT STD_LOGIC;
      in1_rsc_dat : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      in1_rsc_triosy_lz : OUT STD_LOGIC;
      out1_rsc_dat : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
      out1_rsc_triosy_lz : OUT STD_LOGIC;
      coeffs_rsci_radr_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      coeffs_rsci_q_d : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
      coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL fir_core_inst_in1_rsc_dat : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL fir_core_inst_out1_rsc_dat : STD_LOGIC_VECTOR (15 DOWNTO 0);
  SIGNAL fir_core_inst_coeffs_rsci_radr_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL fir_core_inst_coeffs_rsci_q_d : STD_LOGIC_VECTOR (15 DOWNTO 0);

BEGIN
  coeffs_rsci : fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen
    PORT MAP(
      q => coeffs_rsci_q,
      radr => coeffs_rsci_radr,
      radr_d => coeffs_rsci_radr_d_1,
      q_d => coeffs_rsci_q_d_1,
      rport_r_ram_ir_internal_RMASK_B_d => coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d
    );
  coeffs_rsci_q <= coeffs_rsc_q;
  coeffs_rsc_radr <= coeffs_rsci_radr;
  coeffs_rsci_radr_d_1 <= coeffs_rsci_radr_d;
  coeffs_rsci_q_d <= coeffs_rsci_q_d_1;

  fir_core_inst : fir_core
    PORT MAP(
      clk => clk,
      rst => rst,
      coeffs_rsc_triosy_lz => coeffs_rsc_triosy_lz,
      in1_rsc_dat => fir_core_inst_in1_rsc_dat,
      in1_rsc_triosy_lz => in1_rsc_triosy_lz,
      out1_rsc_dat => fir_core_inst_out1_rsc_dat,
      out1_rsc_triosy_lz => out1_rsc_triosy_lz,
      coeffs_rsci_radr_d => fir_core_inst_coeffs_rsci_radr_d,
      coeffs_rsci_q_d => fir_core_inst_coeffs_rsci_q_d,
      coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d => coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d
    );
  fir_core_inst_in1_rsc_dat <= in1_rsc_dat;
  out1_rsc_dat <= fir_core_inst_out1_rsc_dat;
  coeffs_rsci_radr_d <= fir_core_inst_coeffs_rsci_radr_d;
  fir_core_inst_coeffs_rsci_q_d <= coeffs_rsci_q_d;

END v14;



