// nios_system_tb.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module nios_system_tb (
	);

	wire         nios_system_inst_clk_bfm_clk_clk;                   // nios_system_inst_clk_bfm:clk -> [new_sdram_controller_0_my_partner:clk, nios_system_inst:clk_clk, nios_system_inst_reset_bfm:clk]
	wire         nios_system_inst_new_sdram_controller_0_wire_cs_n;  // nios_system_inst:new_sdram_controller_0_wire_cs_n -> new_sdram_controller_0_my_partner:zs_cs_n
	wire   [3:0] nios_system_inst_new_sdram_controller_0_wire_dqm;   // nios_system_inst:new_sdram_controller_0_wire_dqm -> new_sdram_controller_0_my_partner:zs_dqm
	wire         nios_system_inst_new_sdram_controller_0_wire_cas_n; // nios_system_inst:new_sdram_controller_0_wire_cas_n -> new_sdram_controller_0_my_partner:zs_cas_n
	wire         nios_system_inst_new_sdram_controller_0_wire_ras_n; // nios_system_inst:new_sdram_controller_0_wire_ras_n -> new_sdram_controller_0_my_partner:zs_ras_n
	wire         nios_system_inst_new_sdram_controller_0_wire_we_n;  // nios_system_inst:new_sdram_controller_0_wire_we_n -> new_sdram_controller_0_my_partner:zs_we_n
	wire  [12:0] nios_system_inst_new_sdram_controller_0_wire_addr;  // nios_system_inst:new_sdram_controller_0_wire_addr -> new_sdram_controller_0_my_partner:zs_addr
	wire         nios_system_inst_new_sdram_controller_0_wire_cke;   // nios_system_inst:new_sdram_controller_0_wire_cke -> new_sdram_controller_0_my_partner:zs_cke
	wire  [31:0] new_sdram_controller_0_my_partner_conduit_dq;       // [] -> [new_sdram_controller_0_my_partner:zs_dq, nios_system_inst:new_sdram_controller_0_wire_dq]
	wire   [1:0] nios_system_inst_new_sdram_controller_0_wire_ba;    // nios_system_inst:new_sdram_controller_0_wire_ba -> new_sdram_controller_0_my_partner:zs_ba
	wire         nios_system_inst_reset_bfm_reset_reset;             // nios_system_inst_reset_bfm:reset -> nios_system_inst:reset_reset_n

	altera_sdram_partner_module new_sdram_controller_0_my_partner (
		.clk      (nios_system_inst_clk_bfm_clk_clk),                   //     clk.clk
		.zs_dq    (new_sdram_controller_0_my_partner_conduit_dq),       // conduit.dq
		.zs_addr  (nios_system_inst_new_sdram_controller_0_wire_addr),  //        .addr
		.zs_ba    (nios_system_inst_new_sdram_controller_0_wire_ba),    //        .ba
		.zs_cas_n (nios_system_inst_new_sdram_controller_0_wire_cas_n), //        .cas_n
		.zs_cke   (nios_system_inst_new_sdram_controller_0_wire_cke),   //        .cke
		.zs_cs_n  (nios_system_inst_new_sdram_controller_0_wire_cs_n),  //        .cs_n
		.zs_dqm   (nios_system_inst_new_sdram_controller_0_wire_dqm),   //        .dqm
		.zs_ras_n (nios_system_inst_new_sdram_controller_0_wire_ras_n), //        .ras_n
		.zs_we_n  (nios_system_inst_new_sdram_controller_0_wire_we_n)   //        .we_n
	);

	nios_system nios_system_inst (
		.clk_clk                           (nios_system_inst_clk_bfm_clk_clk),                   //                         clk.clk
		.new_sdram_controller_0_wire_addr  (nios_system_inst_new_sdram_controller_0_wire_addr),  // new_sdram_controller_0_wire.addr
		.new_sdram_controller_0_wire_ba    (nios_system_inst_new_sdram_controller_0_wire_ba),    //                            .ba
		.new_sdram_controller_0_wire_cas_n (nios_system_inst_new_sdram_controller_0_wire_cas_n), //                            .cas_n
		.new_sdram_controller_0_wire_cke   (nios_system_inst_new_sdram_controller_0_wire_cke),   //                            .cke
		.new_sdram_controller_0_wire_cs_n  (nios_system_inst_new_sdram_controller_0_wire_cs_n),  //                            .cs_n
		.new_sdram_controller_0_wire_dq    (new_sdram_controller_0_my_partner_conduit_dq),       //                            .dq
		.new_sdram_controller_0_wire_dqm   (nios_system_inst_new_sdram_controller_0_wire_dqm),   //                            .dqm
		.new_sdram_controller_0_wire_ras_n (nios_system_inst_new_sdram_controller_0_wire_ras_n), //                            .ras_n
		.new_sdram_controller_0_wire_we_n  (nios_system_inst_new_sdram_controller_0_wire_we_n),  //                            .we_n
		.reset_reset_n                     (nios_system_inst_reset_bfm_reset_reset),             //                       reset.reset_n
		.sram_0_external_interface_DQ      (),                                                   //   sram_0_external_interface.DQ
		.sram_0_external_interface_ADDR    (),                                                   //                            .ADDR
		.sram_0_external_interface_LB_N    (),                                                   //                            .LB_N
		.sram_0_external_interface_UB_N    (),                                                   //                            .UB_N
		.sram_0_external_interface_CE_N    (),                                                   //                            .CE_N
		.sram_0_external_interface_OE_N    (),                                                   //                            .OE_N
		.sram_0_external_interface_WE_N    ()                                                    //                            .WE_N
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_system_inst_clk_bfm (
		.clk (nios_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nios_system_inst_reset_bfm (
		.reset (nios_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nios_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
