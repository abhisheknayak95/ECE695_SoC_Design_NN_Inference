
//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/mgc_in_wire_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_wire_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule


//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.3d/815731 Production Release
//  HLS Date:       Wed Apr 24 14:54:19 PDT 2019
// 
//  Generated by:   695r48@ecegrid-thin4.ecn.purdue.edu
//  Generated date: Sat Nov 13 22:47:04 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_core_core_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [34:0] fsm_output;
  reg [34:0] fsm_output;


  // FSM State Type Declaration for fir_core_core_fsm_1
  parameter
    main_C_0 = 6'd0,
    main_C_1 = 6'd1,
    main_C_2 = 6'd2,
    main_C_3 = 6'd3,
    main_C_4 = 6'd4,
    main_C_5 = 6'd5,
    main_C_6 = 6'd6,
    main_C_7 = 6'd7,
    main_C_8 = 6'd8,
    main_C_9 = 6'd9,
    main_C_10 = 6'd10,
    main_C_11 = 6'd11,
    main_C_12 = 6'd12,
    main_C_13 = 6'd13,
    main_C_14 = 6'd14,
    main_C_15 = 6'd15,
    main_C_16 = 6'd16,
    main_C_17 = 6'd17,
    main_C_18 = 6'd18,
    main_C_19 = 6'd19,
    main_C_20 = 6'd20,
    main_C_21 = 6'd21,
    main_C_22 = 6'd22,
    main_C_23 = 6'd23,
    main_C_24 = 6'd24,
    main_C_25 = 6'd25,
    main_C_26 = 6'd26,
    main_C_27 = 6'd27,
    main_C_28 = 6'd28,
    main_C_29 = 6'd29,
    main_C_30 = 6'd30,
    main_C_31 = 6'd31,
    main_C_32 = 6'd32,
    main_C_33 = 6'd33,
    main_C_34 = 6'd34;

  reg [5:0] state_var;
  reg [5:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_core_core_fsm_1
    case (state_var)
      main_C_1 : begin
        fsm_output = 35'b00000000000000000000000000000000010;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 35'b00000000000000000000000000000000100;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 35'b00000000000000000000000000000001000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 35'b00000000000000000000000000000010000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 35'b00000000000000000000000000000100000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 35'b00000000000000000000000000001000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 35'b00000000000000000000000000010000000;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 35'b00000000000000000000000000100000000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 35'b00000000000000000000000001000000000;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 35'b00000000000000000000000010000000000;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 35'b00000000000000000000000100000000000;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 35'b00000000000000000000001000000000000;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 35'b00000000000000000000010000000000000;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 35'b00000000000000000000100000000000000;
        state_var_NS = main_C_15;
      end
      main_C_15 : begin
        fsm_output = 35'b00000000000000000001000000000000000;
        state_var_NS = main_C_16;
      end
      main_C_16 : begin
        fsm_output = 35'b00000000000000000010000000000000000;
        state_var_NS = main_C_17;
      end
      main_C_17 : begin
        fsm_output = 35'b00000000000000000100000000000000000;
        state_var_NS = main_C_18;
      end
      main_C_18 : begin
        fsm_output = 35'b00000000000000001000000000000000000;
        state_var_NS = main_C_19;
      end
      main_C_19 : begin
        fsm_output = 35'b00000000000000010000000000000000000;
        state_var_NS = main_C_20;
      end
      main_C_20 : begin
        fsm_output = 35'b00000000000000100000000000000000000;
        state_var_NS = main_C_21;
      end
      main_C_21 : begin
        fsm_output = 35'b00000000000001000000000000000000000;
        state_var_NS = main_C_22;
      end
      main_C_22 : begin
        fsm_output = 35'b00000000000010000000000000000000000;
        state_var_NS = main_C_23;
      end
      main_C_23 : begin
        fsm_output = 35'b00000000000100000000000000000000000;
        state_var_NS = main_C_24;
      end
      main_C_24 : begin
        fsm_output = 35'b00000000001000000000000000000000000;
        state_var_NS = main_C_25;
      end
      main_C_25 : begin
        fsm_output = 35'b00000000010000000000000000000000000;
        state_var_NS = main_C_26;
      end
      main_C_26 : begin
        fsm_output = 35'b00000000100000000000000000000000000;
        state_var_NS = main_C_27;
      end
      main_C_27 : begin
        fsm_output = 35'b00000001000000000000000000000000000;
        state_var_NS = main_C_28;
      end
      main_C_28 : begin
        fsm_output = 35'b00000010000000000000000000000000000;
        state_var_NS = main_C_29;
      end
      main_C_29 : begin
        fsm_output = 35'b00000100000000000000000000000000000;
        state_var_NS = main_C_30;
      end
      main_C_30 : begin
        fsm_output = 35'b00001000000000000000000000000000000;
        state_var_NS = main_C_31;
      end
      main_C_31 : begin
        fsm_output = 35'b00010000000000000000000000000000000;
        state_var_NS = main_C_32;
      end
      main_C_32 : begin
        fsm_output = 35'b00100000000000000000000000000000000;
        state_var_NS = main_C_33;
      end
      main_C_33 : begin
        fsm_output = 35'b01000000000000000000000000000000000;
        state_var_NS = main_C_34;
      end
      main_C_34 : begin
        fsm_output = 35'b10000000000000000000000000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 35'b00000000000000000000000000000000001;
        state_var_NS = main_C_1;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, coeffs_rsc_z, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz, out1_rsc_dat,
      out1_rsc_triosy_lz
);
  input clk;
  input rst;
  input [511:0] coeffs_rsc_z;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;


  // Interconnect Declarations
  wire [511:0] coeffs_rsci_d;
  wire [15:0] in1_rsci_idat;
  reg [15:0] out1_rsci_idat;
  reg out1_rsc_triosy_obj_ld;
  wire [34:0] fsm_output;
  reg [495:0] reg_MAC_io_read_coeffs_rsc_ftd_16;
  reg reg_in1_rsc_triosy_obj_ld_cse;
  reg [15:0] reg_MAC_asn_88_cse;
  reg [15:0] reg_MAC_asn_87_cse;
  reg [15:0] reg_MAC_asn_86_cse;
  reg [15:0] reg_MAC_asn_85_cse;
  reg [15:0] reg_MAC_asn_84_cse;
  reg [15:0] reg_MAC_asn_83_cse;
  reg [15:0] reg_MAC_asn_82_cse;
  reg [15:0] reg_MAC_asn_81_cse;
  reg [15:0] reg_MAC_asn_80_cse;
  reg [15:0] reg_MAC_asn_79_cse;
  reg [15:0] reg_MAC_asn_78_cse;
  reg [15:0] reg_MAC_asn_77_cse;
  reg [15:0] reg_MAC_asn_76_cse;
  reg [15:0] reg_MAC_asn_75_cse;
  reg [15:0] reg_MAC_asn_74_cse;
  reg [15:0] reg_MAC_asn_73_cse;
  reg [15:0] reg_MAC_asn_72_cse;
  reg [15:0] reg_MAC_asn_71_cse;
  reg [15:0] reg_MAC_asn_70_cse;
  reg [15:0] reg_MAC_asn_69_cse;
  reg [15:0] reg_MAC_asn_68_cse;
  reg [15:0] reg_MAC_asn_67_cse;
  reg [15:0] reg_MAC_asn_66_cse;
  reg [15:0] reg_MAC_asn_65_cse;
  reg [15:0] reg_MAC_asn_64_cse;
  reg [15:0] reg_MAC_asn_63_cse;
  reg [15:0] reg_MAC_asn_62_cse;
  wire [29:0] z_out;
  wire [30:0] nl_z_out;
  wire [29:0] z_out_2;
  wire signed [31:0] nl_z_out_2;
  wire [29:0] z_out_3;
  wire signed [31:0] nl_z_out_3;
  reg [15:0] regs_2_sva;
  reg [15:0] regs_30_sva;
  reg [15:0] regs_0_sva;
  reg [29:0] MAC_acc_29_itm;
  reg [29:0] MAC_11_mul_itm;
  reg [29:0] MAC_acc_23_itm;
  reg [29:0] MAC_acc_11_itm;
  reg [15:0] MAC_asn_89_itm;
  reg [15:0] MAC_asn_90_itm;
  reg [29:0] MAC_acc_18_itm;
  wire [30:0] nl_MAC_acc_18_itm;
  wire [29:0] MAC_acc_25_itm_mx0w5;
  wire [30:0] nl_MAC_acc_25_itm_mx0w5;
  wire MAC_acc_11_itm_mx0c5;
  wire MAC_acc_23_itm_mx0c0;
  wire MAC_or_4_cse;

  wire[29:0] mul_nl;
  wire signed [31:0] nl_mul_nl;
  wire[15:0] MAC_mux1h_12_nl;
  wire[0:0] MAC_or_15_nl;
  wire[15:0] MAC_mux1h_13_nl;
  wire[29:0] MAC_acc_16_nl;
  wire[30:0] nl_MAC_acc_16_nl;
  wire[29:0] MAC_4_mul_nl;
  wire signed [31:0] nl_MAC_4_mul_nl;
  wire[29:0] MAC_acc_14_nl;
  wire[30:0] nl_MAC_acc_14_nl;
  wire[29:0] MAC_8_mul_nl;
  wire signed [31:0] nl_MAC_8_mul_nl;
  wire[29:0] mul_3_nl;
  wire signed [31:0] nl_mul_3_nl;
  wire[15:0] MAC_mux1h_16_nl;
  wire[15:0] MAC_mux1h_17_nl;
  wire[29:0] MAC_acc_12_nl;
  wire[30:0] nl_MAC_acc_12_nl;
  wire[29:0] MAC_12_mul_nl;
  wire signed [31:0] nl_MAC_12_mul_nl;
  wire[29:0] MAC_acc_10_nl;
  wire[30:0] nl_MAC_acc_10_nl;
  wire[29:0] MAC_16_mul_nl;
  wire signed [31:0] nl_MAC_16_mul_nl;
  wire[29:0] mul_4_nl;
  wire signed [31:0] nl_mul_4_nl;
  wire[15:0] MAC_mux1h_18_nl;
  wire[15:0] MAC_mux1h_19_nl;
  wire[29:0] MAC_acc_8_nl;
  wire[30:0] nl_MAC_acc_8_nl;
  wire[29:0] MAC_20_mul_nl;
  wire signed [31:0] nl_MAC_20_mul_nl;
  wire[29:0] MAC_acc_6_nl;
  wire[30:0] nl_MAC_acc_6_nl;
  wire[29:0] MAC_24_mul_nl;
  wire signed [31:0] nl_MAC_24_mul_nl;
  wire[29:0] MAC_acc_4_nl;
  wire[30:0] nl_MAC_acc_4_nl;
  wire[29:0] MAC_28_mul_nl;
  wire signed [31:0] nl_MAC_28_mul_nl;
  wire[29:0] MAC_acc_3_nl;
  wire[30:0] nl_MAC_acc_3_nl;
  wire[29:0] MAC_30_mul_nl;
  wire signed [31:0] nl_MAC_30_mul_nl;
  wire[29:0] MAC_acc_nl;
  wire[30:0] nl_MAC_acc_nl;
  wire[29:0] MAC_acc_30_nl;
  wire[30:0] nl_MAC_acc_30_nl;
  wire[29:0] MAC_acc_26_nl;
  wire[30:0] nl_MAC_acc_26_nl;
  wire[0:0] MAC_or_10_nl;
  wire[0:0] MAC_or_11_nl;
  wire[0:0] MAC_or_12_nl;
  wire[0:0] MAC_or_13_nl;
  wire[29:0] MAC_acc_17_nl;
  wire[30:0] nl_MAC_acc_17_nl;
  wire[29:0] MAC_2_mul_nl;
  wire signed [31:0] nl_MAC_2_mul_nl;
  wire[29:0] MAC_acc_15_nl;
  wire[30:0] nl_MAC_acc_15_nl;
  wire[29:0] MAC_6_mul_nl;
  wire signed [31:0] nl_MAC_6_mul_nl;
  wire[29:0] MAC_acc_13_nl;
  wire[30:0] nl_MAC_acc_13_nl;
  wire[29:0] MAC_10_mul_nl;
  wire signed [31:0] nl_MAC_10_mul_nl;
  wire[29:0] MAC_acc_11_nl;
  wire[30:0] nl_MAC_acc_11_nl;
  wire[29:0] MAC_14_mul_nl;
  wire signed [31:0] nl_MAC_14_mul_nl;
  wire[29:0] MAC_acc_9_nl;
  wire[30:0] nl_MAC_acc_9_nl;
  wire[29:0] MAC_18_mul_nl;
  wire signed [31:0] nl_MAC_18_mul_nl;
  wire[29:0] MAC_acc_5_nl;
  wire[30:0] nl_MAC_acc_5_nl;
  wire[29:0] MAC_26_mul_nl;
  wire signed [31:0] nl_MAC_26_mul_nl;
  wire[29:0] MAC_acc_7_nl;
  wire[30:0] nl_MAC_acc_7_nl;
  wire[29:0] MAC_acc_27_nl;
  wire[30:0] nl_MAC_acc_27_nl;
  wire[29:0] MAC_acc_31_nl;
  wire[30:0] nl_MAC_acc_31_nl;
  wire[29:0] MAC_mux_6_nl;
  wire[0:0] MAC_or_14_nl;
  wire[29:0] MAC_mux_7_nl;
  wire[15:0] MAC_mux_8_nl;
  wire[15:0] MAC_mux_9_nl;
  wire[15:0] MAC_mux1h_14_nl;
  wire[15:0] MAC_mux1h_15_nl;

  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_v2 #(.rscid(32'sd1),
  .width(32'sd512)) coeffs_rsci (
      .d(coeffs_rsci_d),
      .z(coeffs_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd16)) in1_rsci (
      .dat(in1_rsc_dat),
      .idat(in1_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd16)) out1_rsci (
      .idat(out1_rsci_idat),
      .dat(out1_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) coeffs_rsc_triosy_obj (
      .ld(reg_in1_rsc_triosy_obj_ld_cse),
      .lz(coeffs_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) in1_rsc_triosy_obj (
      .ld(reg_in1_rsc_triosy_obj_ld_cse),
      .lz(in1_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) out1_rsc_triosy_obj (
      .ld(out1_rsc_triosy_obj_ld),
      .lz(out1_rsc_triosy_lz)
    );
  fir_core_core_fsm fir_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign MAC_or_4_cse = (fsm_output[18]) | (fsm_output[10]);
  assign nl_MAC_acc_25_itm_mx0w5 = MAC_acc_11_itm + MAC_11_mul_itm;
  assign MAC_acc_25_itm_mx0w5 = nl_MAC_acc_25_itm_mx0w5[29:0];
  assign MAC_acc_11_itm_mx0c5 = (fsm_output[30]) | (fsm_output[22]);
  assign MAC_acc_23_itm_mx0c0 = (fsm_output[14]) | (fsm_output[6]);
  always @(posedge clk) begin
    if ( rst ) begin
      out1_rsci_idat <= 16'b0000000000000000;
    end
    else if ( fsm_output[33] ) begin
      out1_rsci_idat <= z_out[29:14];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_88_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_88_cse <= reg_MAC_asn_87_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_87_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_87_cse <= reg_MAC_asn_86_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_86_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_86_cse <= reg_MAC_asn_85_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_85_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_85_cse <= reg_MAC_asn_84_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_84_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_84_cse <= reg_MAC_asn_83_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_83_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_83_cse <= reg_MAC_asn_82_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_82_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_82_cse <= reg_MAC_asn_81_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_81_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_81_cse <= reg_MAC_asn_80_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_80_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_80_cse <= reg_MAC_asn_79_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_79_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_79_cse <= reg_MAC_asn_78_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_78_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_78_cse <= reg_MAC_asn_77_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_77_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_77_cse <= reg_MAC_asn_76_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_76_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_76_cse <= reg_MAC_asn_75_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_75_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_75_cse <= reg_MAC_asn_74_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_74_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_74_cse <= reg_MAC_asn_73_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_73_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_73_cse <= reg_MAC_asn_72_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_72_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_72_cse <= reg_MAC_asn_71_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_71_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_71_cse <= reg_MAC_asn_70_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_70_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_70_cse <= reg_MAC_asn_69_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_69_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_69_cse <= reg_MAC_asn_68_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_68_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_68_cse <= reg_MAC_asn_67_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_67_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_67_cse <= reg_MAC_asn_66_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_66_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_66_cse <= reg_MAC_asn_65_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_65_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_65_cse <= reg_MAC_asn_64_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_64_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_64_cse <= reg_MAC_asn_63_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_63_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_63_cse <= reg_MAC_asn_62_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_asn_62_cse <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      reg_MAC_asn_62_cse <= regs_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_2_sva <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      regs_2_sva <= MAC_asn_89_itm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( fsm_output[2] ) begin
      regs_0_sva <= MAC_asn_90_itm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_asn_89_itm <= 16'b0000000000000000;
    end
    else if ( (fsm_output[34]) | (fsm_output[2]) ) begin
      MAC_asn_89_itm <= MUX_v_16_2_2(regs_0_sva, reg_MAC_asn_88_cse, fsm_output[34]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out1_rsc_triosy_obj_ld <= 1'b0;
      reg_in1_rsc_triosy_obj_ld_cse <= 1'b0;
      MAC_11_mul_itm <= 30'b000000000000000000000000000000;
    end
    else begin
      out1_rsc_triosy_obj_ld <= fsm_output[33];
      reg_in1_rsc_triosy_obj_ld_cse <= fsm_output[0];
      MAC_11_mul_itm <= MUX1HOT_v_30_14_2((mul_nl), z_out_3, (MAC_acc_16_nl), z_out_2,
          (MAC_acc_14_nl), (mul_3_nl), (MAC_acc_12_nl), (MAC_acc_10_nl), (mul_4_nl),
          (MAC_acc_8_nl), (MAC_acc_6_nl), (MAC_acc_4_nl), (MAC_acc_3_nl), (MAC_acc_nl),
          {(MAC_or_10_nl) , (MAC_or_11_nl) , (fsm_output[5]) , (fsm_output[6]) ,
          (fsm_output[9]) , (MAC_or_12_nl) , (fsm_output[13]) , (fsm_output[17])
          , (MAC_or_13_nl) , (fsm_output[21]) , (fsm_output[25]) , (fsm_output[29])
          , (fsm_output[31]) , (fsm_output[32])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_asn_90_itm <= 16'b0000000000000000;
    end
    else if ( (fsm_output[34]) | (fsm_output[0]) ) begin
      MAC_asn_90_itm <= MUX_v_16_2_2(in1_rsci_idat, regs_30_sva, fsm_output[34]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_30_sva <= 16'b0000000000000000;
    end
    else if ( fsm_output[34] ) begin
      regs_30_sva <= reg_MAC_asn_88_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_18_itm <= 30'b000000000000000000000000000000;
    end
    else if ( fsm_output[1] ) begin
      MAC_acc_18_itm <= nl_MAC_acc_18_itm[29:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_11_itm <= 30'b000000000000000000000000000000;
    end
    else if ( (fsm_output[27]) | (fsm_output[19]) | (fsm_output[15]) | (fsm_output[11])
        | (fsm_output[7]) | (fsm_output[3]) | MAC_acc_11_itm_mx0c5 ) begin
      MAC_acc_11_itm <= MUX1HOT_v_30_7_2((MAC_acc_17_nl), (MAC_acc_15_nl), (MAC_acc_13_nl),
          (MAC_acc_11_nl), (MAC_acc_9_nl), MAC_acc_25_itm_mx0w5, (MAC_acc_5_nl),
          {(fsm_output[3]) , (fsm_output[7]) , (fsm_output[11]) , (fsm_output[15])
          , (fsm_output[19]) , MAC_acc_11_itm_mx0c5 , (fsm_output[27])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_23_itm <= 30'b000000000000000000000000000000;
    end
    else if ( (fsm_output[26]) | MAC_acc_23_itm_mx0c0 | (fsm_output[23]) ) begin
      MAC_acc_23_itm <= MUX1HOT_v_30_3_2(MAC_acc_25_itm_mx0w5, (MAC_acc_7_nl), (MAC_acc_27_nl),
          {MAC_acc_23_itm_mx0c0 , (fsm_output[23]) , (fsm_output[26])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_29_itm <= 30'b000000000000000000000000000000;
    end
    else if ( MAC_or_4_cse ) begin
      MAC_acc_29_itm <= MUX_v_30_2_2(z_out, (MAC_acc_31_nl), fsm_output[18]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_io_read_coeffs_rsc_ftd_16 <= 496'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( fsm_output[0] ) begin
      reg_MAC_io_read_coeffs_rsc_ftd_16 <= coeffs_rsci_d[495:0];
    end
  end
  assign MAC_or_15_nl = (fsm_output[0]) | (fsm_output[2]);
  assign MAC_mux1h_12_nl = MUX1HOT_v_16_3_2(MAC_asn_90_itm, reg_MAC_asn_65_cse, reg_MAC_asn_67_cse,
      {(MAC_or_15_nl) , (fsm_output[8]) , (fsm_output[10])});
  assign MAC_mux1h_13_nl = MUX1HOT_v_16_4_2((coeffs_rsci_d[511:496]), (reg_MAC_io_read_coeffs_rsc_ftd_16[15:0]),
      (reg_MAC_io_read_coeffs_rsc_ftd_16[111:96]), (reg_MAC_io_read_coeffs_rsc_ftd_16[143:128]),
      {(fsm_output[0]) , (fsm_output[2]) , (fsm_output[8]) , (fsm_output[10])});
  assign nl_mul_nl = $signed((MAC_mux1h_12_nl)) * $signed((MAC_mux1h_13_nl));
  assign mul_nl = nl_mul_nl[29:0];
  assign nl_MAC_4_mul_nl = $signed(reg_MAC_asn_62_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[63:48]));
  assign MAC_4_mul_nl = nl_MAC_4_mul_nl[29:0];
  assign nl_MAC_acc_16_nl = MAC_11_mul_itm + (MAC_4_mul_nl);
  assign MAC_acc_16_nl = nl_MAC_acc_16_nl[29:0];
  assign nl_MAC_8_mul_nl = $signed(reg_MAC_asn_66_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[127:112]));
  assign MAC_8_mul_nl = nl_MAC_8_mul_nl[29:0];
  assign nl_MAC_acc_14_nl = MAC_11_mul_itm + (MAC_8_mul_nl);
  assign MAC_acc_14_nl = nl_MAC_acc_14_nl[29:0];
  assign MAC_mux1h_16_nl = MUX1HOT_v_16_4_2(reg_MAC_asn_69_cse, reg_MAC_asn_71_cse,
      reg_MAC_asn_73_cse, reg_MAC_asn_75_cse, {(fsm_output[12]) , (fsm_output[14])
      , (fsm_output[16]) , (fsm_output[18])});
  assign MAC_mux1h_17_nl = MUX1HOT_v_16_4_2((reg_MAC_io_read_coeffs_rsc_ftd_16[175:160]),
      (reg_MAC_io_read_coeffs_rsc_ftd_16[207:192]), (reg_MAC_io_read_coeffs_rsc_ftd_16[239:224]),
      (reg_MAC_io_read_coeffs_rsc_ftd_16[271:256]), {(fsm_output[12]) , (fsm_output[14])
      , (fsm_output[16]) , (fsm_output[18])});
  assign nl_mul_3_nl = $signed((MAC_mux1h_16_nl)) * $signed((MAC_mux1h_17_nl));
  assign mul_3_nl = nl_mul_3_nl[29:0];
  assign nl_MAC_12_mul_nl = $signed(reg_MAC_asn_70_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[191:176]));
  assign MAC_12_mul_nl = nl_MAC_12_mul_nl[29:0];
  assign nl_MAC_acc_12_nl = MAC_11_mul_itm + (MAC_12_mul_nl);
  assign MAC_acc_12_nl = nl_MAC_acc_12_nl[29:0];
  assign nl_MAC_16_mul_nl = $signed(reg_MAC_asn_74_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[255:240]));
  assign MAC_16_mul_nl = nl_MAC_16_mul_nl[29:0];
  assign nl_MAC_acc_10_nl = MAC_11_mul_itm + (MAC_16_mul_nl);
  assign MAC_acc_10_nl = nl_MAC_acc_10_nl[29:0];
  assign MAC_mux1h_18_nl = MUX1HOT_v_16_4_2(reg_MAC_asn_77_cse, reg_MAC_asn_79_cse,
      reg_MAC_asn_81_cse, reg_MAC_asn_83_cse, {(fsm_output[20]) , (fsm_output[22])
      , (fsm_output[24]) , (fsm_output[26])});
  assign MAC_mux1h_19_nl = MUX1HOT_v_16_4_2((reg_MAC_io_read_coeffs_rsc_ftd_16[303:288]),
      (reg_MAC_io_read_coeffs_rsc_ftd_16[335:320]), (reg_MAC_io_read_coeffs_rsc_ftd_16[367:352]),
      (reg_MAC_io_read_coeffs_rsc_ftd_16[399:384]), {(fsm_output[20]) , (fsm_output[22])
      , (fsm_output[24]) , (fsm_output[26])});
  assign nl_mul_4_nl = $signed((MAC_mux1h_18_nl)) * $signed((MAC_mux1h_19_nl));
  assign mul_4_nl = nl_mul_4_nl[29:0];
  assign nl_MAC_20_mul_nl = $signed(reg_MAC_asn_78_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[319:304]));
  assign MAC_20_mul_nl = nl_MAC_20_mul_nl[29:0];
  assign nl_MAC_acc_8_nl = MAC_11_mul_itm + (MAC_20_mul_nl);
  assign MAC_acc_8_nl = nl_MAC_acc_8_nl[29:0];
  assign nl_MAC_24_mul_nl = $signed(reg_MAC_asn_82_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[383:368]));
  assign MAC_24_mul_nl = nl_MAC_24_mul_nl[29:0];
  assign nl_MAC_acc_6_nl = MAC_11_mul_itm + (MAC_24_mul_nl);
  assign MAC_acc_6_nl = nl_MAC_acc_6_nl[29:0];
  assign nl_MAC_28_mul_nl = $signed(reg_MAC_asn_86_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[447:432]));
  assign MAC_28_mul_nl = nl_MAC_28_mul_nl[29:0];
  assign nl_MAC_acc_4_nl = MAC_11_mul_itm + (MAC_28_mul_nl);
  assign MAC_acc_4_nl = nl_MAC_acc_4_nl[29:0];
  assign nl_MAC_30_mul_nl = $signed(reg_MAC_asn_88_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[479:464]));
  assign MAC_30_mul_nl = nl_MAC_30_mul_nl[29:0];
  assign nl_MAC_acc_3_nl = MAC_11_mul_itm + (MAC_30_mul_nl);
  assign MAC_acc_3_nl = nl_MAC_acc_3_nl[29:0];
  assign nl_MAC_acc_26_nl = MAC_11_mul_itm + MAC_acc_18_itm;
  assign MAC_acc_26_nl = nl_MAC_acc_26_nl[29:0];
  assign nl_MAC_acc_30_nl = MAC_acc_11_itm + (MAC_acc_26_nl);
  assign MAC_acc_30_nl = nl_MAC_acc_30_nl[29:0];
  assign nl_MAC_acc_nl = MAC_acc_23_itm + (MAC_acc_30_nl);
  assign MAC_acc_nl = nl_MAC_acc_nl[29:0];
  assign MAC_or_10_nl = (fsm_output[0]) | (fsm_output[2]) | (fsm_output[8]) | (fsm_output[10]);
  assign MAC_or_11_nl = (fsm_output[4]) | (fsm_output[28]) | (fsm_output[30]);
  assign MAC_or_12_nl = (fsm_output[12]) | (fsm_output[14]) | (fsm_output[16]) |
      (fsm_output[18]);
  assign MAC_or_13_nl = (fsm_output[20]) | (fsm_output[22]) | (fsm_output[24]) |
      (fsm_output[26]);
  assign nl_MAC_acc_18_itm  = z_out_3 + MAC_11_mul_itm;
  assign nl_MAC_2_mul_nl = $signed(MAC_asn_89_itm) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[31:16]));
  assign MAC_2_mul_nl = nl_MAC_2_mul_nl[29:0];
  assign nl_MAC_acc_17_nl = MAC_11_mul_itm + (MAC_2_mul_nl);
  assign MAC_acc_17_nl = nl_MAC_acc_17_nl[29:0];
  assign nl_MAC_6_mul_nl = $signed(reg_MAC_asn_64_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[95:80]));
  assign MAC_6_mul_nl = nl_MAC_6_mul_nl[29:0];
  assign nl_MAC_acc_15_nl = MAC_11_mul_itm + (MAC_6_mul_nl);
  assign MAC_acc_15_nl = nl_MAC_acc_15_nl[29:0];
  assign nl_MAC_10_mul_nl = $signed(reg_MAC_asn_68_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[159:144]));
  assign MAC_10_mul_nl = nl_MAC_10_mul_nl[29:0];
  assign nl_MAC_acc_13_nl = MAC_11_mul_itm + (MAC_10_mul_nl);
  assign MAC_acc_13_nl = nl_MAC_acc_13_nl[29:0];
  assign nl_MAC_14_mul_nl = $signed(reg_MAC_asn_72_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[223:208]));
  assign MAC_14_mul_nl = nl_MAC_14_mul_nl[29:0];
  assign nl_MAC_acc_11_nl = MAC_11_mul_itm + (MAC_14_mul_nl);
  assign MAC_acc_11_nl = nl_MAC_acc_11_nl[29:0];
  assign nl_MAC_18_mul_nl = $signed(reg_MAC_asn_76_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[287:272]));
  assign MAC_18_mul_nl = nl_MAC_18_mul_nl[29:0];
  assign nl_MAC_acc_9_nl = MAC_11_mul_itm + (MAC_18_mul_nl);
  assign MAC_acc_9_nl = nl_MAC_acc_9_nl[29:0];
  assign nl_MAC_26_mul_nl = $signed(reg_MAC_asn_84_cse) * $signed((reg_MAC_io_read_coeffs_rsc_ftd_16[415:400]));
  assign MAC_26_mul_nl = nl_MAC_26_mul_nl[29:0];
  assign nl_MAC_acc_5_nl = MAC_11_mul_itm + (MAC_26_mul_nl);
  assign MAC_acc_5_nl = nl_MAC_acc_5_nl[29:0];
  assign nl_MAC_acc_7_nl = MAC_11_mul_itm + z_out_2;
  assign MAC_acc_7_nl = nl_MAC_acc_7_nl[29:0];
  assign nl_MAC_acc_27_nl = MAC_acc_11_itm + z_out;
  assign MAC_acc_27_nl = nl_MAC_acc_27_nl[29:0];
  assign nl_MAC_acc_31_nl = MAC_acc_29_itm + z_out;
  assign MAC_acc_31_nl = nl_MAC_acc_31_nl[29:0];
  assign MAC_or_14_nl = (fsm_output[26]) | MAC_or_4_cse;
  assign MAC_mux_6_nl = MUX_v_30_2_2(MAC_acc_29_itm, MAC_acc_23_itm, MAC_or_14_nl);
  assign MAC_mux_7_nl = MUX_v_30_2_2(MAC_11_mul_itm, MAC_acc_25_itm_mx0w5, MAC_or_4_cse);
  assign nl_z_out = (MAC_mux_6_nl) + (MAC_mux_7_nl);
  assign z_out = nl_z_out[29:0];
  assign MAC_mux_8_nl = MUX_v_16_2_2(reg_MAC_asn_63_cse, reg_MAC_asn_80_cse, fsm_output[23]);
  assign MAC_mux_9_nl = MUX_v_16_2_2((reg_MAC_io_read_coeffs_rsc_ftd_16[79:64]),
      (reg_MAC_io_read_coeffs_rsc_ftd_16[351:336]), fsm_output[23]);
  assign nl_z_out_2 = $signed((MAC_mux_8_nl)) * $signed((MAC_mux_9_nl));
  assign z_out_2 = nl_z_out_2[29:0];
  assign MAC_mux1h_14_nl = MUX1HOT_v_16_4_2(regs_2_sva, reg_MAC_asn_85_cse, reg_MAC_asn_87_cse,
      MAC_asn_89_itm, {(fsm_output[4]) , (fsm_output[28]) , (fsm_output[30]) , (fsm_output[1])});
  assign MAC_mux1h_15_nl = MUX1HOT_v_16_4_2((reg_MAC_io_read_coeffs_rsc_ftd_16[47:32]),
      (reg_MAC_io_read_coeffs_rsc_ftd_16[431:416]), (reg_MAC_io_read_coeffs_rsc_ftd_16[463:448]),
      (reg_MAC_io_read_coeffs_rsc_ftd_16[495:480]), {(fsm_output[4]) , (fsm_output[28])
      , (fsm_output[30]) , (fsm_output[1])});
  assign nl_z_out_3 = $signed((MAC_mux1h_14_nl)) * $signed((MAC_mux1h_15_nl));
  assign z_out_3 = nl_z_out_3[29:0];

  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_4_2;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [3:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    MUX1HOT_v_16_4_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_14_2;
    input [29:0] input_13;
    input [29:0] input_12;
    input [29:0] input_11;
    input [29:0] input_10;
    input [29:0] input_9;
    input [29:0] input_8;
    input [29:0] input_7;
    input [29:0] input_6;
    input [29:0] input_5;
    input [29:0] input_4;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [13:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    result = result | ( input_3 & {30{sel[3]}});
    result = result | ( input_4 & {30{sel[4]}});
    result = result | ( input_5 & {30{sel[5]}});
    result = result | ( input_6 & {30{sel[6]}});
    result = result | ( input_7 & {30{sel[7]}});
    result = result | ( input_8 & {30{sel[8]}});
    result = result | ( input_9 & {30{sel[9]}});
    result = result | ( input_10 & {30{sel[10]}});
    result = result | ( input_11 & {30{sel[11]}});
    result = result | ( input_12 & {30{sel[12]}});
    result = result | ( input_13 & {30{sel[13]}});
    MUX1HOT_v_30_14_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_3_2;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [2:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    MUX1HOT_v_30_3_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_7_2;
    input [29:0] input_6;
    input [29:0] input_5;
    input [29:0] input_4;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [6:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    result = result | ( input_3 & {30{sel[3]}});
    result = result | ( input_4 & {30{sel[4]}});
    result = result | ( input_5 & {30{sel[5]}});
    result = result | ( input_6 & {30{sel[6]}});
    MUX1HOT_v_30_7_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, coeffs_rsc_z, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz, out1_rsc_dat,
      out1_rsc_triosy_lz
);
  input clk;
  input rst;
  input [511:0] coeffs_rsc_z;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .coeffs_rsc_z(coeffs_rsc_z),
      .coeffs_rsc_triosy_lz(coeffs_rsc_triosy_lz),
      .in1_rsc_dat(in1_rsc_dat),
      .in1_rsc_triosy_lz(in1_rsc_triosy_lz),
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_triosy_lz(out1_rsc_triosy_lz)
    );
endmodule



