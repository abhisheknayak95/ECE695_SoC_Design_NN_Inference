
//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.3d/815731 Production Release
//  HLS Date:       Wed Apr 24 14:54:19 PDT 2019
// 
//  Generated by:   695r48@cparch23.ecn.purdue.edu
//  Generated date: Tue Nov  9 15:18:43 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen
// ------------------------------------------------------------------


module fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen (
  q, radr, radr_d, q_d, rport_r_ram_ir_internal_RMASK_B_d
);
  input [15:0] q;
  output [4:0] radr;
  input [4:0] radr_d;
  output [15:0] q_d;
  input rport_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_core_core_fsm (
  clk, rst, fsm_output, MAC_C_3_tr0
);
  input clk;
  input rst;
  output [19:0] fsm_output;
  reg [19:0] fsm_output;
  input MAC_C_3_tr0;


  // FSM State Type Declaration for fir_core_core_fsm_1
  parameter
    main_C_0 = 5'd0,
    MAC_C_0 = 5'd1,
    MAC_C_1 = 5'd2,
    MAC_C_2 = 5'd3,
    MAC_C_3 = 5'd4,
    MAC_C_4 = 5'd5,
    MAC_C_5 = 5'd6,
    MAC_C_6 = 5'd7,
    MAC_C_7 = 5'd8,
    MAC_C_8 = 5'd9,
    MAC_C_9 = 5'd10,
    MAC_C_10 = 5'd11,
    MAC_C_11 = 5'd12,
    MAC_C_12 = 5'd13,
    MAC_C_13 = 5'd14,
    MAC_C_14 = 5'd15,
    MAC_C_15 = 5'd16,
    MAC_C_16 = 5'd17,
    MAC_C_17 = 5'd18,
    main_C_1 = 5'd19;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_core_core_fsm_1
    case (state_var)
      MAC_C_0 : begin
        fsm_output = 20'b00000000000000000010;
        state_var_NS = MAC_C_1;
      end
      MAC_C_1 : begin
        fsm_output = 20'b00000000000000000100;
        state_var_NS = MAC_C_2;
      end
      MAC_C_2 : begin
        fsm_output = 20'b00000000000000001000;
        state_var_NS = MAC_C_3;
      end
      MAC_C_3 : begin
        fsm_output = 20'b00000000000000010000;
        if ( MAC_C_3_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = MAC_C_4;
        end
      end
      MAC_C_4 : begin
        fsm_output = 20'b00000000000000100000;
        state_var_NS = MAC_C_5;
      end
      MAC_C_5 : begin
        fsm_output = 20'b00000000000001000000;
        state_var_NS = MAC_C_6;
      end
      MAC_C_6 : begin
        fsm_output = 20'b00000000000010000000;
        state_var_NS = MAC_C_7;
      end
      MAC_C_7 : begin
        fsm_output = 20'b00000000000100000000;
        state_var_NS = MAC_C_8;
      end
      MAC_C_8 : begin
        fsm_output = 20'b00000000001000000000;
        state_var_NS = MAC_C_9;
      end
      MAC_C_9 : begin
        fsm_output = 20'b00000000010000000000;
        state_var_NS = MAC_C_10;
      end
      MAC_C_10 : begin
        fsm_output = 20'b00000000100000000000;
        state_var_NS = MAC_C_11;
      end
      MAC_C_11 : begin
        fsm_output = 20'b00000001000000000000;
        state_var_NS = MAC_C_12;
      end
      MAC_C_12 : begin
        fsm_output = 20'b00000010000000000000;
        state_var_NS = MAC_C_13;
      end
      MAC_C_13 : begin
        fsm_output = 20'b00000100000000000000;
        state_var_NS = MAC_C_14;
      end
      MAC_C_14 : begin
        fsm_output = 20'b00001000000000000000;
        state_var_NS = MAC_C_15;
      end
      MAC_C_15 : begin
        fsm_output = 20'b00010000000000000000;
        state_var_NS = MAC_C_16;
      end
      MAC_C_16 : begin
        fsm_output = 20'b00100000000000000000;
        state_var_NS = MAC_C_17;
      end
      MAC_C_17 : begin
        fsm_output = 20'b01000000000000000000;
        state_var_NS = MAC_C_0;
      end
      main_C_1 : begin
        fsm_output = 20'b10000000000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 20'b00000000000000000001;
        state_var_NS = MAC_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz, out1_rsc_dat, out1_rsc_triosy_lz,
      coeffs_rsci_radr_d, coeffs_rsci_q_d, coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d
);
  input clk;
  input rst;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;
  output [4:0] coeffs_rsci_radr_d;
  input [15:0] coeffs_rsci_q_d;
  output coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire [15:0] in1_rsci_idat;
  reg [15:0] out1_rsci_idat;
  wire [19:0] fsm_output;
  wire [5:0] MAC_2_acc_2_tmp;
  wire [6:0] nl_MAC_2_acc_2_tmp;
  wire or_dcpl_1;
  wire and_dcpl_4;
  wire and_dcpl_21;
  wire and_dcpl_22;
  wire and_dcpl_24;
  wire and_dcpl_31;
  wire and_dcpl_36;
  wire or_dcpl_45;
  wire or_dcpl_56;
  wire or_dcpl_61;
  wire or_dcpl_62;
  wire or_dcpl_63;
  wire or_dcpl_67;
  wire and_dcpl_39;
  wire or_tmp_178;
  wire or_tmp_183;
  wire or_tmp_197;
  wire or_tmp_199;
  wire [1:0] MAC_acc_7_psp_1_sva_1;
  wire [2:0] nl_MAC_acc_7_psp_1_sva_1;
  wire [2:0] MAC_acc_3_psp_sva_1;
  wire [3:0] nl_MAC_acc_3_psp_sva_1;
  wire MAC_i_or_cse;
  reg reg_out1_rsc_triosy_obj_ld_cse;
  wire reg_out1_out1_and_cse;
  reg [1:0] MAC_acc_10_psp_sva;
  wire [4:0] MAC_1_acc_2_psp_sva_mx0w0;
  wire [5:0] nl_MAC_1_acc_2_psp_sva_mx0w0;
  reg MAC_i_4_0_sva_4;
  reg MAC_i_4_0_sva_0;
  reg [3:0] MAC_acc_psp_sva;
  wire [4:0] nl_MAC_acc_psp_sva;
  reg [2:0] MAC_acc_9_psp_sva;
  reg [2:0] MAC_acc_3_psp_sva;
  reg [1:0] MAC_acc_4_psp_sva;
  reg [1:0] MAC_acc_7_psp_1_sva;
  wire [29:0] z_out;
  wire [30:0] nl_z_out;
  wire [29:0] z_out_1;
  wire [30:0] nl_z_out_1;
  wire [15:0] z_out_2;
  wire [29:0] z_out_4;
  wire signed [31:0] nl_z_out_4;
  wire [29:0] z_out_5;
  wire signed [31:0] nl_z_out_5;
  wire [29:0] z_out_6;
  wire signed [31:0] nl_z_out_6;
  wire [29:0] z_out_7;
  wire signed [31:0] nl_z_out_7;
  wire [4:0] z_out_9;
  wire [5:0] nl_z_out_9;
  reg [15:0] regs_15_sva;
  reg [15:0] regs_16_sva;
  reg [15:0] regs_14_sva;
  reg [15:0] regs_17_sva;
  reg [15:0] regs_13_sva;
  reg [15:0] regs_18_sva;
  reg [15:0] regs_12_sva;
  reg [15:0] regs_19_sva;
  reg [15:0] regs_11_sva;
  reg [15:0] regs_20_sva;
  reg [15:0] regs_10_sva;
  reg [15:0] regs_21_sva;
  reg [15:0] regs_9_sva;
  reg [15:0] regs_22_sva;
  reg [15:0] regs_8_sva;
  reg [15:0] regs_23_sva;
  reg [15:0] regs_7_sva;
  reg [15:0] regs_24_sva;
  reg [15:0] regs_6_sva;
  reg [15:0] regs_25_sva;
  reg [15:0] regs_5_sva;
  reg [15:0] regs_26_sva;
  reg [15:0] regs_4_sva;
  reg [15:0] regs_27_sva;
  reg [15:0] regs_3_sva;
  reg [15:0] regs_28_sva;
  reg [15:0] regs_2_sva;
  reg [15:0] regs_29_sva;
  reg [15:0] regs_1_sva;
  reg [15:0] regs_30_sva;
  reg [15:0] regs_0_sva;
  reg [29:0] acc_32_3_1_sva;
  reg [15:0] regs_30_sva_1;
  reg [15:0] regs_29_sva_1;
  reg [15:0] regs_28_sva_1;
  reg [15:0] regs_27_sva_1;
  reg [15:0] regs_26_sva_1;
  reg [15:0] regs_25_sva_1;
  reg [15:0] regs_24_sva_1;
  reg [15:0] regs_23_sva_1;
  reg [15:0] regs_22_sva_1;
  reg [15:0] regs_21_sva_1;
  reg [15:0] regs_20_sva_1;
  reg [15:0] regs_19_sva_1;
  reg [15:0] regs_18_sva_1;
  reg [15:0] regs_17_sva_1;
  reg [15:0] regs_16_sva_1;
  reg [15:0] regs_15_sva_1;
  reg [15:0] regs_14_sva_1;
  reg [15:0] regs_13_sva_1;
  reg [15:0] regs_12_sva_1;
  reg [15:0] regs_11_sva_1;
  reg [15:0] regs_10_sva_1;
  reg [15:0] regs_9_sva_1;
  reg [15:0] regs_8_sva_1;
  reg [15:0] regs_7_sva_1;
  reg [15:0] regs_6_sva_1;
  reg [15:0] regs_5_sva_1;
  reg [15:0] regs_4_sva_1;
  reg [15:0] regs_3_sva_1;
  reg [15:0] regs_2_sva_1;
  reg [15:0] regs_1_sva_1;
  reg [15:0] regs_0_sva_1;
  reg [15:0] MAC_4_MAC_mux_itm;
  reg [29:0] MAC_4_mul_itm;
  reg [15:0] MAC_5_MAC_mux_itm;
  reg [15:0] MAC_6_MAC_mux_itm;
  reg [15:0] MAC_7_MAC_mux_itm;
  reg [15:0] MAC_8_MAC_mux_itm;
  reg [15:0] MAC_mux_2_itm;
  reg [15:0] MAC_10_MAC_mux_itm;
  reg [29:0] MAC_10_mul_itm;
  reg [15:0] MAC_11_MAC_mux_itm;
  reg [29:0] MAC_11_mul_itm;
  reg [29:0] MAC_acc_14_itm;
  reg [29:0] MAC_acc_20_itm;
  reg [15:0] MAC_12_MAC_mux_itm;
  reg [15:0] MAC_13_MAC_mux_itm;
  reg [15:0] MAC_14_MAC_mux_itm;
  reg [15:0] MAC_15_MAC_mux_itm;
  reg [15:0] MAC_3_MAC_mux_itm;
  reg [29:0] MAC_acc_18_itm;
  wire [30:0] nl_MAC_acc_18_itm;
  wire [29:0] MAC_acc_11_mx0w2;
  wire [30:0] nl_MAC_acc_11_mx0w2;
  wire [4:0] MAC_9_acc_2_psp_sva_1;
  wire [5:0] nl_MAC_9_acc_2_psp_sva_1;
  wire [1:0] MAC_acc_4_psp_sva_1;
  wire [2:0] nl_MAC_acc_4_psp_sva_1;
  wire [2:0] MAC_acc_9_psp_sva_1;
  wire [3:0] nl_MAC_acc_9_psp_sva_1;
  wire or_281_tmp;
  wire or_276_tmp;
  wire nor_16_tmp;
  wire or_262_tmp;
  wire and_480_tmp;
  reg reg_MAC_15_acc_2_ftd;
  reg reg_MAC_15_acc_2_ftd_4;
  wire MAC_and_20_rgt;
  wire MAC_and_21_rgt;
  wire MAC_and_22_rgt;
  wire MAC_and_23_rgt;
  wire MAC_and_14_rgt;
  wire MAC_and_15_rgt;
  wire MAC_and_16_rgt;
  wire MAC_and_17_rgt;
  reg [1:0] MAC_i_5_0_3_sva_rsp_0;
  reg [1:0] MAC_i_5_0_3_sva_rsp_2;
  reg MAC_13_acc_2_psp_sva_rsp_0;
  reg MAC_13_acc_2_psp_sva_rsp_2;
  wire reg_MAC_13_acc_2_psp_rgt_ssc;
  reg MAC_9_acc_2_psp_sva_rsp_0;
  reg MAC_9_acc_2_psp_sva_rsp_2;
  wire MAC_and_m1c;
  wire MAC_and_m1c_1;
  wire MAC_and_m1c_2;
  wire MAC_conc_146_tmp_2;
  wire [1:0] MAC_conc_146_tmp_1_0;

  wire[29:0] acc_mux1h_1_nl;
  wire[0:0] acc_not_nl;
  wire[0:0] MAC_MAC_or_nl;
  wire[1:0] MAC_acc_10_nl;
  wire[2:0] nl_MAC_acc_10_nl;
  wire[0:0] MAC_and_42_nl;
  wire[0:0] MAC_and_40_nl;
  wire[0:0] MAC_and_35_nl;
  wire[0:0] MAC_and_36_nl;
  wire[0:0] MAC_and_37_nl;
  wire[0:0] MAC_and_38_nl;
  wire[0:0] MAC_and_34_nl;
  wire[0:0] MAC_MAC_nor_7_nl;
  wire[0:0] MAC_and_29_nl;
  wire[0:0] MAC_and_3_nl;
  wire[0:0] MAC_and_4_nl;
  wire[0:0] MAC_and_5_nl;
  wire[0:0] MAC_and_24_nl;
  wire[0:0] MAC_and_25_nl;
  wire[0:0] MAC_and_26_nl;
  wire[0:0] MAC_and_27_nl;
  wire[0:0] MAC_and_nl;
  wire[0:0] MAC_and_1_nl;
  wire[0:0] MAC_and_2_nl;
  wire[0:0] MAC_and_19_nl;
  wire[0:0] MAC_and_10_nl;
  wire[0:0] MAC_and_11_nl;
  wire[0:0] MAC_and_12_nl;
  wire[0:0] MAC_and_13_nl;
  wire[29:0] mul_nl;
  wire signed [31:0] nl_mul_nl;
  wire[15:0] MAC_mux_46_nl;
  wire[29:0] MAC_acc_22_nl;
  wire[30:0] nl_MAC_acc_22_nl;
  wire[29:0] MAC_acc_19_nl;
  wire[30:0] nl_MAC_acc_19_nl;
  wire[0:0] MAC_or_nl;
  wire[0:0] MAC_or_12_nl;
  wire[0:0] MAC_or_13_nl;
  wire[29:0] mul_5_nl;
  wire signed [31:0] nl_mul_5_nl;
  wire[15:0] MAC_mux_51_nl;
  wire[29:0] MAC_8_mul_nl;
  wire signed [31:0] nl_MAC_8_mul_nl;
  wire[0:0] MAC_or_10_nl;
  wire[29:0] MAC_acc_23_nl;
  wire[30:0] nl_MAC_acc_23_nl;
  wire[29:0] MAC_acc_21_nl;
  wire[30:0] nl_MAC_acc_21_nl;
  wire[0:0] MAC_mux1h_3_nl;
  wire[0:0] MAC_or_2_nl;
  wire[0:0] MAC_or_3_nl;
  wire[0:0] MAC_or_7_nl;
  wire[0:0] MAC_or_4_nl;
  wire[0:0] MAC_mux1h_54_nl;
  wire[0:0] MAC_or_5_nl;
  wire[0:0] MAC_mux1h_56_nl;
  wire[0:0] MAC_or_6_nl;
  wire[0:0] MAC_mux1h_57_nl;
  wire[0:0] MAC_mux1h_55_nl;
  wire[29:0] MAC_mux_45_nl;
  wire[15:0] MAC_mux_47_nl;
  wire[0:0] or_326_nl;
  wire[15:0] MAC_mux_48_nl;
  wire[0:0] or_327_nl;
  wire[15:0] MAC_mux_49_nl;
  wire[15:0] MAC_mux_50_nl;
  wire[0:0] MAC_mux_52_nl;
  wire[0:0] MAC_MAC_or_2_nl;
  wire[1:0] MAC_mux_53_nl;
  wire[0:0] MAC_and_43_nl;
  wire[0:0] MAC_and_44_nl;
  wire[0:0] MAC_and_45_nl;
  wire[0:0] MAC_and_46_nl;
  wire[0:0] MAC_and_47_nl;
  wire[0:0] MAC_and_48_nl;
  wire[0:0] MAC_and_49_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_fir_core_core_fsm_inst_MAC_C_3_tr0;
  assign nl_fir_core_core_fsm_inst_MAC_C_3_tr0 = MAC_i_5_0_3_sva_rsp_0[1];
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd16)) in1_rsci (
      .dat(in1_rsc_dat),
      .idat(in1_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd16)) out1_rsci (
      .idat(out1_rsci_idat),
      .dat(out1_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) coeffs_rsc_triosy_obj (
      .ld(reg_out1_rsc_triosy_obj_ld_cse),
      .lz(coeffs_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) in1_rsc_triosy_obj (
      .ld(reg_out1_rsc_triosy_obj_ld_cse),
      .lz(in1_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) out1_rsc_triosy_obj (
      .ld(reg_out1_rsc_triosy_obj_ld_cse),
      .lz(out1_rsc_triosy_lz)
    );
  fir_core_core_fsm fir_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .MAC_C_3_tr0(nl_fir_core_core_fsm_inst_MAC_C_3_tr0[0:0])
    );
  assign reg_out1_out1_and_cse = (fsm_output[4]) & (MAC_i_5_0_3_sva_rsp_0[1]);
  assign MAC_i_or_cse = (fsm_output[0]) | (fsm_output[4]);
  assign MAC_and_20_rgt = ~((z_out_9[4]) | (z_out_9[0]) | nor_16_tmp);
  assign MAC_and_21_rgt = (z_out_9[0]) & (~ (z_out_9[4])) & (~ nor_16_tmp);
  assign MAC_and_22_rgt = (z_out_9[4]) & (~ (z_out_9[0])) & (~ nor_16_tmp);
  assign MAC_and_23_rgt = (z_out_9[4]) & (z_out_9[0]) & (~ nor_16_tmp);
  assign MAC_and_14_rgt = ~((MAC_9_acc_2_psp_sva_1[4]) | (~ (MAC_acc_4_psp_sva_1[0]))
      | or_tmp_199);
  assign MAC_and_15_rgt = ~((MAC_acc_4_psp_sva_1[0]) | (MAC_9_acc_2_psp_sva_1[4])
      | or_tmp_199);
  assign MAC_and_16_rgt = (MAC_9_acc_2_psp_sva_1[4]) & (MAC_acc_4_psp_sva_1[0]) &
      (~ or_tmp_199);
  assign MAC_and_17_rgt = (MAC_9_acc_2_psp_sva_1[4]) & (~ (MAC_acc_4_psp_sva_1[0]))
      & (~ or_tmp_199);
  assign nl_MAC_acc_11_mx0w2 = MAC_10_mul_itm + MAC_11_mul_itm;
  assign MAC_acc_11_mx0w2 = nl_MAC_acc_11_mx0w2[29:0];
  assign nl_MAC_1_acc_2_psp_sva_mx0w0 = ({MAC_i_4_0_sva_4 , (signext_3_1(MAC_acc_10_psp_sva[0]))
      , MAC_i_4_0_sva_0}) + 5'b00001;
  assign MAC_1_acc_2_psp_sva_mx0w0 = nl_MAC_1_acc_2_psp_sva_mx0w0[4:0];
  assign nl_MAC_2_acc_2_tmp = conv_u2s_5_6(MAC_1_acc_2_psp_sva_mx0w0) + 6'b000001;
  assign MAC_2_acc_2_tmp = nl_MAC_2_acc_2_tmp[5:0];
  assign nl_MAC_acc_3_psp_sva_1 = conv_u2u_2_3({1'b1 , (~ (MAC_2_acc_2_tmp[0]))})
      + 3'b001;
  assign MAC_acc_3_psp_sva_1 = nl_MAC_acc_3_psp_sva_1[2:0];
  assign nl_MAC_acc_7_psp_1_sva_1 = conv_u2u_1_2(~ (MAC_acc_3_psp_sva_1[0])) + 2'b01;
  assign MAC_acc_7_psp_1_sva_1 = nl_MAC_acc_7_psp_1_sva_1[1:0];
  assign nl_MAC_9_acc_2_psp_sva_1 = ({(MAC_i_5_0_3_sva_rsp_0[0]) , MAC_acc_psp_sva})
      + 5'b00001;
  assign MAC_9_acc_2_psp_sva_1 = nl_MAC_9_acc_2_psp_sva_1[4:0];
  assign nl_MAC_acc_4_psp_sva_1 = conv_u2u_1_2(MAC_9_acc_2_psp_sva_1[0]) + 2'b01;
  assign MAC_acc_4_psp_sva_1 = nl_MAC_acc_4_psp_sva_1[1:0];
  assign nl_MAC_acc_9_psp_sva_1 = conv_u2u_2_3({1'b1 , (~ (MAC_acc_4_psp_sva_1[0]))})
      + 3'b001;
  assign MAC_acc_9_psp_sva_1 = nl_MAC_acc_9_psp_sva_1[2:0];
  assign or_dcpl_1 = (fsm_output[7:6]!=2'b00);
  assign and_dcpl_4 = ~((fsm_output[19]) | (fsm_output[0]));
  assign and_dcpl_21 = ~((fsm_output[18:17]!=2'b00));
  assign and_dcpl_22 = and_dcpl_21 & (~ (fsm_output[16]));
  assign and_dcpl_24 = ~((fsm_output[2:1]!=2'b00));
  assign and_dcpl_31 = ~((fsm_output[0]) | (fsm_output[14]) | (fsm_output[15]) |
      (fsm_output[1]));
  assign and_dcpl_36 = and_dcpl_21 & (~ (fsm_output[16])) & (~ (fsm_output[19]));
  assign or_dcpl_45 = (fsm_output[4:3]!=2'b00);
  assign or_dcpl_56 = (fsm_output[8:7]!=2'b00);
  assign or_dcpl_61 = (fsm_output[3:2]!=2'b00);
  assign or_dcpl_62 = or_dcpl_61 | (fsm_output[4]);
  assign or_dcpl_63 = (fsm_output[5]) | (fsm_output[8]);
  assign or_dcpl_67 = (fsm_output[6]) | (fsm_output[3]) | (fsm_output[4]);
  assign and_dcpl_39 = ~((fsm_output[0]) | (fsm_output[15]));
  assign or_tmp_178 = and_dcpl_22 & (~ (fsm_output[19])) & (~ (fsm_output[13])) &
      and_dcpl_31;
  assign or_tmp_183 = (fsm_output[5]) | (fsm_output[10]) | (fsm_output[9]) | or_dcpl_56
      | (fsm_output[6]) | (fsm_output[2]) | or_dcpl_45;
  assign or_tmp_197 = (fsm_output[7:5]!=3'b000) | or_dcpl_45;
  assign or_tmp_199 = (fsm_output[6:5]!=2'b00) | or_dcpl_45;
  assign MAC_or_2_nl = (fsm_output[3]) | (fsm_output[9]) | (fsm_output[10]) | (fsm_output[11])
      | (fsm_output[12]) | (fsm_output[13]);
  assign MAC_or_3_nl = (fsm_output[8:5]!=4'b0000);
  assign MAC_or_7_nl = (fsm_output[15:14]!=2'b00);
  assign MAC_mux1h_3_nl = MUX1HOT_s_1_6_2((MAC_1_acc_2_psp_sva_mx0w0[4]), MAC_i_4_0_sva_4,
      (MAC_i_5_0_3_sva_rsp_0[0]), (MAC_i_5_0_3_sva_rsp_0[0]), MAC_9_acc_2_psp_sva_rsp_0,
      MAC_13_acc_2_psp_sva_rsp_0, {(fsm_output[1]) , (fsm_output[2]) , (MAC_or_2_nl)
      , (fsm_output[4]) , (MAC_or_3_nl) , (MAC_or_7_nl)});
  assign MAC_mux1h_54_nl = MUX1HOT_s_1_3_2((MAC_1_acc_2_psp_sva_mx0w0[3]), (MAC_acc_10_psp_sva[0]),
      (MAC_acc_psp_sva[3]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[9])});
  assign MAC_or_4_nl = ((MAC_mux1h_54_nl) & (~ (fsm_output[4])) & (~((fsm_output[3])
      | (fsm_output[10]) | (fsm_output[11]) | (fsm_output[12]) | (fsm_output[13]))))
      | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[14])
      | (fsm_output[15]);
  assign MAC_mux1h_56_nl = MUX1HOT_s_1_5_2((MAC_1_acc_2_psp_sva_mx0w0[2]), (MAC_acc_10_psp_sva[0]),
      (MAC_acc_9_psp_sva[2]), (MAC_acc_psp_sva[2]), (MAC_acc_3_psp_sva[2]), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[9]) , (fsm_output[13])});
  assign MAC_or_5_nl = ((MAC_mux1h_56_nl) & (~ (fsm_output[4])) & (~((fsm_output[3])
      | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8])))) | (fsm_output[10])
      | (fsm_output[11]) | (fsm_output[12]) | (fsm_output[14]) | (fsm_output[15]);
  assign MAC_mux1h_57_nl = MUX1HOT_s_1_9_2((MAC_1_acc_2_psp_sva_mx0w0[1]), (MAC_acc_10_psp_sva[0]),
      (MAC_i_5_0_3_sva_rsp_2[1]), (MAC_acc_9_psp_sva[1]), (MAC_acc_4_psp_sva[1]),
      (MAC_acc_psp_sva[1]), (MAC_acc_7_psp_1_sva[1]), (MAC_acc_3_psp_sva[1]), (MAC_acc_10_psp_sva[1]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13]) , (fsm_output[14])});
  assign MAC_or_6_nl = ((MAC_mux1h_57_nl) & (~((fsm_output[8]) | (fsm_output[12])
      | (fsm_output[15])))) | (fsm_output[3]) | (fsm_output[6]) | (fsm_output[10]);
  assign MAC_mux1h_55_nl = MUX1HOT_s_1_15_2((MAC_1_acc_2_psp_sva_mx0w0[0]), MAC_i_4_0_sva_0,
      (~ (MAC_i_5_0_3_sva_rsp_2[0])), (MAC_i_5_0_3_sva_rsp_2[0]), (MAC_acc_9_psp_sva[0]),
      (~ (MAC_acc_4_psp_sva[0])), (MAC_acc_4_psp_sva[0]), MAC_9_acc_2_psp_sva_rsp_2,
      (MAC_acc_psp_sva[0]), (~ (MAC_acc_7_psp_1_sva[0])), (MAC_acc_7_psp_1_sva[0]),
      (~ (MAC_acc_3_psp_sva[0])), (MAC_acc_3_psp_sva[0]), (MAC_acc_10_psp_sva[0]),
      MAC_13_acc_2_psp_sva_rsp_2, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])
      , (fsm_output[9]) , (fsm_output[10]) , (fsm_output[11]) , (fsm_output[12])
      , (fsm_output[13]) , (fsm_output[14]) , (fsm_output[15])});
  assign coeffs_rsci_radr_d = {(MAC_mux1h_3_nl) , (MAC_or_4_nl) , (MAC_or_5_nl) ,
      (MAC_or_6_nl) , (MAC_mux1h_55_nl)};
  assign coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d = (and_dcpl_22 & and_dcpl_4
      & (~ (fsm_output[4]))) | ((~ (MAC_i_5_0_3_sva_rsp_0[1])) & (fsm_output[4]));
  assign and_480_tmp = and_dcpl_36 & and_dcpl_31;
  assign or_262_tmp = (fsm_output[11]) | (fsm_output[5]) | (fsm_output[10]) | (fsm_output[9])
      | (fsm_output[8]) | or_dcpl_1 | (fsm_output[2]) | or_dcpl_45;
  assign nor_16_tmp = ~((~ and_dcpl_36) | (fsm_output[2:0]!=3'b000));
  assign reg_MAC_13_acc_2_psp_rgt_ssc = ~(and_dcpl_36 & and_dcpl_39 & and_dcpl_24);
  assign or_276_tmp = (fsm_output[5]) | (fsm_output[9]) | or_dcpl_56 | or_dcpl_67;
  assign or_281_tmp = (fsm_output[5:3]!=3'b000);
  always @(posedge clk) begin
    if ( rst ) begin
      acc_32_3_1_sva <= 30'b000000000000000000000000000000;
    end
    else if ( (fsm_output[18]) | (fsm_output[0]) | (fsm_output[8]) | (fsm_output[4])
        ) begin
      acc_32_3_1_sva <= MUX_v_30_2_2(30'b000000000000000000000000000000, (acc_mux1h_1_nl),
          (acc_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out1_rsci_idat <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
      regs_15_sva <= 16'b0000000000000000;
      regs_30_sva <= 16'b0000000000000000;
      regs_14_sva <= 16'b0000000000000000;
      regs_29_sva <= 16'b0000000000000000;
      regs_13_sva <= 16'b0000000000000000;
      regs_28_sva <= 16'b0000000000000000;
      regs_11_sva <= 16'b0000000000000000;
      regs_12_sva <= 16'b0000000000000000;
      regs_27_sva <= 16'b0000000000000000;
      regs_10_sva <= 16'b0000000000000000;
      regs_26_sva <= 16'b0000000000000000;
      regs_9_sva <= 16'b0000000000000000;
      regs_25_sva <= 16'b0000000000000000;
      regs_8_sva <= 16'b0000000000000000;
      regs_24_sva <= 16'b0000000000000000;
      regs_7_sva <= 16'b0000000000000000;
      regs_23_sva <= 16'b0000000000000000;
      regs_22_sva <= 16'b0000000000000000;
      regs_16_sva <= 16'b0000000000000000;
      regs_1_sva <= 16'b0000000000000000;
      regs_6_sva <= 16'b0000000000000000;
      regs_21_sva <= 16'b0000000000000000;
      regs_4_sva <= 16'b0000000000000000;
      regs_5_sva <= 16'b0000000000000000;
      regs_20_sva <= 16'b0000000000000000;
      regs_19_sva <= 16'b0000000000000000;
      regs_18_sva <= 16'b0000000000000000;
      regs_3_sva <= 16'b0000000000000000;
      regs_2_sva <= 16'b0000000000000000;
      regs_17_sva <= 16'b0000000000000000;
    end
    else if ( reg_out1_out1_and_cse ) begin
      out1_rsci_idat <= z_out_1[29:14];
      regs_0_sva <= regs_0_sva_1;
      regs_15_sva <= regs_15_sva_1;
      regs_30_sva <= regs_30_sva_1;
      regs_14_sva <= regs_14_sva_1;
      regs_29_sva <= regs_29_sva_1;
      regs_13_sva <= regs_13_sva_1;
      regs_28_sva <= regs_28_sva_1;
      regs_11_sva <= regs_11_sva_1;
      regs_12_sva <= regs_12_sva_1;
      regs_27_sva <= regs_27_sva_1;
      regs_10_sva <= regs_10_sva_1;
      regs_26_sva <= regs_26_sva_1;
      regs_9_sva <= regs_9_sva_1;
      regs_25_sva <= regs_25_sva_1;
      regs_8_sva <= regs_8_sva_1;
      regs_24_sva <= regs_24_sva_1;
      regs_7_sva <= regs_7_sva_1;
      regs_23_sva <= regs_23_sva_1;
      regs_22_sva <= regs_22_sva_1;
      regs_16_sva <= regs_16_sva_1;
      regs_1_sva <= regs_1_sva_1;
      regs_6_sva <= regs_6_sva_1;
      regs_21_sva <= regs_21_sva_1;
      regs_4_sva <= regs_4_sva_1;
      regs_5_sva <= regs_5_sva_1;
      regs_20_sva <= regs_20_sva_1;
      regs_19_sva <= regs_19_sva_1;
      regs_18_sva <= regs_18_sva_1;
      regs_3_sva <= regs_3_sva_1;
      regs_2_sva <= regs_2_sva_1;
      regs_17_sva <= regs_17_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_i_4_0_sva_4 <= 1'b0;
      MAC_i_4_0_sva_0 <= 1'b0;
    end
    else if ( MAC_i_or_cse ) begin
      MAC_i_4_0_sva_4 <= reg_MAC_15_acc_2_ftd & (fsm_output[4]);
      MAC_i_4_0_sva_0 <= reg_MAC_15_acc_2_ftd_4 & (fsm_output[4]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_0_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_0_sva_1 <= in1_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_out1_rsc_triosy_obj_ld_cse <= 1'b0;
      MAC_10_mul_itm <= 30'b000000000000000000000000000000;
    end
    else begin
      reg_out1_rsc_triosy_obj_ld_cse <= reg_out1_out1_and_cse;
      MAC_10_mul_itm <= MUX1HOT_v_30_5_2(z_out_4, (mul_5_nl), z_out_5, (MAC_8_mul_nl),
          z_out_7, {(fsm_output[3]) , (MAC_or_10_nl) , (fsm_output[9]) , (fsm_output[11])
          , (fsm_output[16])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_30_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_30_sva_1 <= regs_29_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_29_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_29_sva_1 <= regs_28_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_28_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_28_sva_1 <= regs_27_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_27_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_27_sva_1 <= regs_26_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_26_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_26_sva_1 <= regs_25_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_25_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_25_sva_1 <= regs_24_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_24_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_24_sva_1 <= regs_23_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_23_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_23_sva_1 <= regs_22_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_22_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_22_sva_1 <= regs_21_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_21_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_21_sva_1 <= regs_20_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_20_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_20_sva_1 <= regs_19_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_19_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_19_sva_1 <= regs_18_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_18_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_18_sva_1 <= regs_17_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_17_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_17_sva_1 <= regs_16_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_16_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_16_sva_1 <= regs_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_15_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_15_sva_1 <= regs_14_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_14_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_14_sva_1 <= regs_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_13_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_13_sva_1 <= regs_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_12_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_12_sva_1 <= regs_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_11_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_11_sva_1 <= regs_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_10_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_10_sva_1 <= regs_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_9_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_9_sva_1 <= regs_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_8_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_8_sva_1 <= regs_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_7_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_7_sva_1 <= regs_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_6_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_6_sva_1 <= regs_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_5_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_5_sva_1 <= regs_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_4_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_4_sva_1 <= regs_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_3_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_3_sva_1 <= regs_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_2_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_2_sva_1 <= regs_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_1_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ and_dcpl_4 ) begin
      regs_1_sva_1 <= regs_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_10_psp_sva <= 2'b00;
    end
    else if ( ~(and_dcpl_22 & and_dcpl_4 & (fsm_output[15:14]==2'b00) & and_dcpl_24)
        ) begin
      MAC_acc_10_psp_sva <= MUX_v_2_2_2(({1'b0 , (MAC_MAC_or_nl)}), (MAC_acc_10_nl),
          fsm_output[2]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_5_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ and_480_tmp ) begin
      MAC_5_MAC_mux_itm <= MUX_v_16_2_2(regs_18_sva, regs_3_sva, MAC_and_42_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_6_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_tmp_178 ) begin
      MAC_6_MAC_mux_itm <= MUX_v_16_2_2(regs_4_sva, regs_19_sva, MAC_and_40_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_3_psp_sva <= 3'b000;
    end
    else if ( ~ or_tmp_178 ) begin
      MAC_acc_3_psp_sva <= MAC_acc_3_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_7_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_262_tmp ) begin
      MAC_7_MAC_mux_itm <= MUX1HOT_v_16_4_2(regs_4_sva, regs_5_sva, regs_20_sva,
          regs_21_sva, {(MAC_and_35_nl) , (MAC_and_36_nl) , (MAC_and_37_nl) , (MAC_and_38_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_tmp_183 ) begin
      MAC_8_MAC_mux_itm <= MUX_v_16_2_2(regs_6_sva, regs_21_sva, MAC_and_34_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_7_psp_1_sva <= 2'b00;
    end
    else if ( ~ or_tmp_183 ) begin
      MAC_acc_7_psp_1_sva <= MAC_acc_7_psp_1_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_psp_sva <= 4'b0000;
    end
    else if ( ~(or_dcpl_63 | or_dcpl_1 | or_dcpl_62) ) begin
      MAC_acc_psp_sva <= nl_MAC_acc_psp_sva[3:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_3_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_62 ) begin
      MAC_3_MAC_mux_itm <= MUX1HOT_v_16_3_2(regs_15_sva, regs_16_sva, regs_1_sva,
          {(MAC_MAC_nor_7_nl) , (MAC_2_acc_2_tmp[0]) , (MAC_2_acc_2_tmp[1])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_4_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_61 ) begin
      MAC_4_MAC_mux_itm <= MUX_v_16_2_2(regs_2_sva, regs_17_sva, MAC_and_29_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_10_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~(or_dcpl_63 | (fsm_output[7]) | or_dcpl_67) ) begin
      MAC_10_MAC_mux_itm <= MUX1HOT_v_16_7_2(regs_0_sva, regs_15_sva, regs_30_sva,
          regs_7_sva, regs_8_sva, regs_23_sva, regs_24_sva, {(MAC_and_3_nl) , (MAC_and_4_nl)
          , (MAC_and_5_nl) , (MAC_and_24_nl) , (MAC_and_25_nl) , (MAC_and_26_nl)
          , (MAC_and_27_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_15_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( (~(and_dcpl_36 & and_dcpl_39 & (~ (fsm_output[1])))) | (fsm_output[3])
        ) begin
      MAC_15_MAC_mux_itm <= MUX1HOT_v_16_4_2(regs_0_sva_1, regs_14_sva, regs_29_sva,
          z_out_2, {(MAC_and_nl) , (MAC_and_1_nl) , (MAC_and_2_nl) , (fsm_output[3])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( MAC_and_20_rgt | MAC_and_21_rgt | MAC_and_22_rgt | MAC_and_23_rgt )
        begin
      MAC_14_MAC_mux_itm <= MUX1HOT_v_16_4_2(regs_11_sva, regs_12_sva, regs_27_sva,
          regs_28_sva, {MAC_and_20_rgt , MAC_and_21_rgt , MAC_and_22_rgt , MAC_and_23_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_mux_2_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_276_tmp ) begin
      MAC_mux_2_itm <= MUX_v_16_2_2(regs_22_sva, regs_7_sva, MAC_and_19_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_11_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_tmp_197 ) begin
      MAC_11_MAC_mux_itm <= z_out_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_12_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( MAC_and_14_rgt | MAC_and_15_rgt | MAC_and_16_rgt | MAC_and_17_rgt )
        begin
      MAC_12_MAC_mux_itm <= MUX1HOT_v_16_4_2(regs_9_sva, regs_10_sva, regs_25_sva,
          regs_26_sva, {MAC_and_14_rgt , MAC_and_15_rgt , MAC_and_16_rgt , MAC_and_17_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_4_psp_sva <= 2'b00;
    end
    else if ( ~ or_tmp_199 ) begin
      MAC_acc_4_psp_sva <= MAC_acc_4_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_13_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_281_tmp ) begin
      MAC_13_MAC_mux_itm <= MUX1HOT_v_16_4_2(regs_10_sva, regs_11_sva, regs_26_sva,
          regs_27_sva, {(MAC_and_10_nl) , (MAC_and_11_nl) , (MAC_and_12_nl) , (MAC_and_13_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_9_psp_sva <= 3'b000;
    end
    else if ( ~ or_dcpl_45 ) begin
      MAC_acc_9_psp_sva <= MAC_acc_9_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_11_mul_itm <= 30'b000000000000000000000000000000;
    end
    else if ( (fsm_output[17]) | (fsm_output[5]) | (fsm_output[12]) | (fsm_output[10])
        | (fsm_output[8]) | (fsm_output[6]) | (fsm_output[2]) | (fsm_output[14])
        | (fsm_output[15]) ) begin
      MAC_11_mul_itm <= MUX1HOT_v_30_6_2(z_out_5, (mul_nl), z_out_4, z_out_6, z_out_7,
          (MAC_acc_22_nl), {(MAC_or_nl) , (MAC_or_12_nl) , (MAC_or_13_nl) , (fsm_output[12])
          , (fsm_output[14]) , (fsm_output[17])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_4_mul_itm <= 30'b000000000000000000000000000000;
    end
    else if ( (fsm_output[15]) | (fsm_output[4]) ) begin
      MAC_4_mul_itm <= MUX_v_30_2_2(z_out_6, (MAC_acc_23_nl), fsm_output[15]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_18_itm <= 30'b000000000000000000000000000000;
    end
    else if ( fsm_output[6] ) begin
      MAC_acc_18_itm <= nl_MAC_acc_18_itm[29:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_14_itm <= 30'b000000000000000000000000000000;
    end
    else if ( (fsm_output[14]) | (fsm_output[10]) ) begin
      MAC_acc_14_itm <= MAC_acc_11_mx0w2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_20_itm <= 30'b000000000000000000000000000000;
    end
    else if ( fsm_output[12] ) begin
      MAC_acc_20_itm <= z_out_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_i_5_0_3_sva_rsp_0 <= 2'b00;
    end
    else if ( ~ or_tmp_178 ) begin
      MAC_i_5_0_3_sva_rsp_0 <= MAC_2_acc_2_tmp[5:4];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_i_5_0_3_sva_rsp_2 <= 2'b00;
    end
    else if ( ~ or_tmp_178 ) begin
      MAC_i_5_0_3_sva_rsp_2 <= MAC_2_acc_2_tmp[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_13_acc_2_psp_sva_rsp_0 <= 1'b0;
      MAC_13_acc_2_psp_sva_rsp_2 <= 1'b0;
    end
    else if ( reg_MAC_13_acc_2_psp_rgt_ssc ) begin
      MAC_13_acc_2_psp_sva_rsp_0 <= z_out_9[4];
      MAC_13_acc_2_psp_sva_rsp_2 <= z_out_9[0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_9_acc_2_psp_sva_rsp_0 <= 1'b0;
    end
    else if ( ~ or_tmp_197 ) begin
      MAC_9_acc_2_psp_sva_rsp_0 <= MAC_9_acc_2_psp_sva_1[4];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_9_acc_2_psp_sva_rsp_2 <= 1'b0;
    end
    else if ( ~ or_tmp_197 ) begin
      MAC_9_acc_2_psp_sva_rsp_2 <= MAC_9_acc_2_psp_sva_1[0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_15_acc_2_ftd <= 1'b0;
    end
    else if ( ~ (MAC_i_5_0_3_sva_rsp_0[1]) ) begin
      reg_MAC_15_acc_2_ftd <= z_out_9[4];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_MAC_15_acc_2_ftd_4 <= 1'b0;
    end
    else if ( ~ (MAC_i_5_0_3_sva_rsp_0[1]) ) begin
      reg_MAC_15_acc_2_ftd_4 <= z_out_9[0];
    end
  end
  assign acc_mux1h_1_nl = MUX1HOT_v_30_3_2(z_out_1, MAC_acc_11_mx0w2, z_out, {(fsm_output[4])
      , (fsm_output[8]) , (fsm_output[18])});
  assign acc_not_nl = ~ (fsm_output[0]);
  assign MAC_mux_51_nl = MUX_v_16_2_2(MAC_12_MAC_mux_itm, MAC_6_MAC_mux_itm, fsm_output[13]);
  assign nl_mul_5_nl = $signed((MAC_mux_51_nl)) * $signed((coeffs_rsci_q_d));
  assign mul_5_nl = nl_mul_5_nl[29:0];
  assign nl_MAC_8_mul_nl = $signed(MAC_8_MAC_mux_itm) * $signed((coeffs_rsci_q_d));
  assign MAC_8_mul_nl = nl_MAC_8_mul_nl[29:0];
  assign MAC_or_10_nl = (fsm_output[7]) | (fsm_output[13]);
  assign MAC_MAC_or_nl = ((MAC_acc_10_psp_sva[0]) & (fsm_output[1])) | (fsm_output[18]);
  assign nl_MAC_acc_10_nl = conv_u2u_1_2(z_out_9[0]) + 2'b01;
  assign MAC_acc_10_nl = nl_MAC_acc_10_nl[1:0];
  assign MAC_and_42_nl = (MAC_acc_3_psp_sva_1==3'b100) & (~ and_480_tmp);
  assign MAC_and_40_nl = (MAC_acc_3_psp_sva_1[0]) & (~ or_tmp_178);
  assign MAC_and_35_nl = (MAC_acc_7_psp_1_sva_1[0]) & (~((MAC_2_acc_2_tmp[4]) | (MAC_acc_7_psp_1_sva_1[1])))
      & (~ or_262_tmp);
  assign MAC_and_36_nl = (MAC_acc_7_psp_1_sva_1[1]) & (~((MAC_2_acc_2_tmp[4]) | (MAC_acc_7_psp_1_sva_1[0])))
      & (~ or_262_tmp);
  assign MAC_and_37_nl = (MAC_2_acc_2_tmp[4]) & (MAC_acc_7_psp_1_sva_1==2'b01) &
      (~ or_262_tmp);
  assign MAC_and_38_nl = (MAC_2_acc_2_tmp[4]) & (MAC_acc_7_psp_1_sva_1==2'b10) &
      (~ or_262_tmp);
  assign MAC_and_34_nl = (MAC_acc_7_psp_1_sva_1[0]) & (~ or_tmp_183);
  assign nl_MAC_acc_psp_sva  = conv_u2u_3_4({2'b11 , (~ (MAC_acc_7_psp_1_sva_1[0]))})
      + 4'b0001;
  assign MAC_MAC_nor_7_nl = ~((MAC_2_acc_2_tmp[1:0]!=2'b00) | or_dcpl_62);
  assign MAC_and_29_nl = (MAC_2_acc_2_tmp[0]) & (~ or_dcpl_61);
  assign MAC_and_3_nl = (MAC_1_acc_2_psp_sva_mx0w0==5'b00001) & (fsm_output[1]);
  assign MAC_and_4_nl = (MAC_1_acc_2_psp_sva_mx0w0==5'b10000) & (fsm_output[1]);
  assign MAC_and_5_nl = (MAC_1_acc_2_psp_sva_mx0w0==5'b11111) & (fsm_output[1]);
  assign MAC_and_24_nl = (~((MAC_9_acc_2_psp_sva_1[4]) | (MAC_9_acc_2_psp_sva_1[0])))
      & (fsm_output[2]);
  assign MAC_and_25_nl = (MAC_9_acc_2_psp_sva_1[0]) & (~ (MAC_9_acc_2_psp_sva_1[4]))
      & (fsm_output[2]);
  assign MAC_and_26_nl = (MAC_9_acc_2_psp_sva_1[4]) & (~ (MAC_9_acc_2_psp_sva_1[0]))
      & (fsm_output[2]);
  assign MAC_and_27_nl = (MAC_9_acc_2_psp_sva_1[4]) & (MAC_9_acc_2_psp_sva_1[0])
      & (fsm_output[2]);
  assign MAC_and_nl = (~(MAC_i_4_0_sva_4 | (MAC_acc_10_psp_sva[0]) | MAC_i_4_0_sva_0))
      & (fsm_output[1]);
  assign MAC_and_1_nl = (MAC_acc_10_psp_sva[0]) & MAC_i_4_0_sva_0 & (~ MAC_i_4_0_sva_4)
      & (fsm_output[1]);
  assign MAC_and_2_nl = MAC_i_4_0_sva_4 & (MAC_acc_10_psp_sva[0]) & (~ MAC_i_4_0_sva_0)
      & (fsm_output[1]);
  assign MAC_and_19_nl = (MAC_acc_psp_sva==4'b1000) & (~ or_276_tmp);
  assign MAC_and_10_nl = (MAC_acc_9_psp_sva_1[1:0]==2'b11) & (~((MAC_9_acc_2_psp_sva_1[4])
      | (MAC_acc_9_psp_sva_1[2]))) & (~ or_281_tmp);
  assign MAC_and_11_nl = (MAC_acc_9_psp_sva_1[2]) & (~((MAC_9_acc_2_psp_sva_1[4])
      | (MAC_acc_9_psp_sva_1[1:0]!=2'b00))) & (~ or_281_tmp);
  assign MAC_and_12_nl = (MAC_9_acc_2_psp_sva_1[4]) & (MAC_acc_9_psp_sva_1==3'b011)
      & (~ or_281_tmp);
  assign MAC_and_13_nl = (MAC_9_acc_2_psp_sva_1[4]) & (MAC_acc_9_psp_sva_1==3'b100)
      & (~ or_281_tmp);
  assign MAC_mux_46_nl = MUX_v_16_2_2(MAC_3_MAC_mux_itm, MAC_13_MAC_mux_itm, fsm_output[6]);
  assign nl_mul_nl = $signed((MAC_mux_46_nl)) * $signed((coeffs_rsci_q_d));
  assign mul_nl = nl_mul_nl[29:0];
  assign nl_MAC_acc_19_nl = acc_32_3_1_sva + MAC_acc_11_mx0w2;
  assign MAC_acc_19_nl = nl_MAC_acc_19_nl[29:0];
  assign nl_MAC_acc_22_nl = (MAC_acc_19_nl) + MAC_acc_18_itm;
  assign MAC_acc_22_nl = nl_MAC_acc_22_nl[29:0];
  assign MAC_or_nl = (fsm_output[2]) | (fsm_output[10]);
  assign MAC_or_12_nl = (fsm_output[6:5]!=2'b00);
  assign MAC_or_13_nl = (fsm_output[8]) | (fsm_output[15]);
  assign nl_MAC_acc_21_nl = z_out + MAC_acc_14_itm;
  assign MAC_acc_21_nl = nl_MAC_acc_21_nl[29:0];
  assign nl_MAC_acc_23_nl = (MAC_acc_21_nl) + MAC_acc_20_itm;
  assign MAC_acc_23_nl = nl_MAC_acc_23_nl[29:0];
  assign nl_MAC_acc_18_itm  = acc_32_3_1_sva + MAC_11_mul_itm;
  assign nl_z_out = MAC_4_mul_itm + MAC_11_mul_itm;
  assign z_out = nl_z_out[29:0];
  assign MAC_mux_45_nl = MUX_v_30_2_2(MAC_acc_14_itm, acc_32_3_1_sva, fsm_output[4]);
  assign nl_z_out_1 = MAC_acc_11_mx0w2 + (MAC_mux_45_nl);
  assign z_out_1 = nl_z_out_1[29:0];
  assign or_326_nl = (fsm_output[15]) | (fsm_output[3]);
  assign MAC_mux_47_nl = MUX_v_16_2_2(MAC_11_MAC_mux_itm, MAC_15_MAC_mux_itm, or_326_nl);
  assign nl_z_out_4 = $signed((MAC_mux_47_nl)) * $signed((coeffs_rsci_q_d));
  assign z_out_4 = nl_z_out_4[29:0];
  assign or_327_nl = (fsm_output[2]) | (fsm_output[9]);
  assign MAC_mux_48_nl = MUX_v_16_2_2(MAC_mux_2_itm, MAC_10_MAC_mux_itm, or_327_nl);
  assign nl_z_out_5 = $signed((MAC_mux_48_nl)) * $signed((coeffs_rsci_q_d));
  assign z_out_5 = nl_z_out_5[29:0];
  assign MAC_mux_49_nl = MUX_v_16_2_2(MAC_7_MAC_mux_itm, MAC_4_MAC_mux_itm, fsm_output[4]);
  assign nl_z_out_6 = $signed((MAC_mux_49_nl)) * $signed((coeffs_rsci_q_d));
  assign z_out_6 = nl_z_out_6[29:0];
  assign MAC_mux_50_nl = MUX_v_16_2_2(MAC_5_MAC_mux_itm, MAC_14_MAC_mux_itm, fsm_output[16]);
  assign nl_z_out_7 = $signed((MAC_mux_50_nl)) * $signed((coeffs_rsci_q_d));
  assign z_out_7 = nl_z_out_7[29:0];
  assign MAC_mux_52_nl = MUX_s_1_2_2((MAC_9_acc_2_psp_sva_1[4]), MAC_13_acc_2_psp_sva_rsp_0,
      fsm_output[3]);
  assign MAC_MAC_or_2_nl = (MAC_acc_9_psp_sva_1[2]) | (fsm_output[3]);
  assign MAC_mux_53_nl = MUX_v_2_2_2((signext_2_1(MAC_acc_9_psp_sva_1[0])), MAC_acc_10_psp_sva,
      fsm_output[3]);
  assign nl_z_out_9 = ({(MAC_mux_52_nl) , 1'b1 , (MAC_MAC_or_2_nl) , (MAC_mux_53_nl)})
      + 5'b00001;
  assign z_out_9 = nl_z_out_9[4:0];
  assign MAC_conc_146_tmp_2 = MUX_s_1_2_2(MAC_13_acc_2_psp_sva_rsp_0, (MAC_9_acc_2_psp_sva_1[4]),
      fsm_output[2]);
  assign MAC_conc_146_tmp_1_0 = MUX_v_2_2_2(MAC_acc_10_psp_sva, MAC_acc_4_psp_sva_1,
      fsm_output[2]);
  assign MAC_and_m1c = (MAC_conc_146_tmp_1_0[1]) & (~(MAC_conc_146_tmp_2 | (MAC_conc_146_tmp_1_0[0])));
  assign MAC_and_m1c_1 = MAC_conc_146_tmp_2 & (MAC_conc_146_tmp_1_0==2'b01);
  assign MAC_and_m1c_2 = MAC_conc_146_tmp_2 & (MAC_conc_146_tmp_1_0==2'b10);
  assign MAC_and_43_nl = (MAC_conc_146_tmp_1_0[0]) & (~(MAC_conc_146_tmp_2 | (MAC_conc_146_tmp_1_0[1])));
  assign MAC_and_44_nl = (~ (fsm_output[2])) & MAC_and_m1c;
  assign MAC_and_45_nl = (fsm_output[2]) & MAC_and_m1c;
  assign MAC_and_46_nl = (~ (fsm_output[2])) & MAC_and_m1c_1;
  assign MAC_and_47_nl = (fsm_output[2]) & MAC_and_m1c_1;
  assign MAC_and_48_nl = (~ (fsm_output[2])) & MAC_and_m1c_2;
  assign MAC_and_49_nl = (fsm_output[2]) & MAC_and_m1c_2;
  assign z_out_2 = MUX1HOT_v_16_7_2(regs_8_sva, regs_13_sva, regs_9_sva, regs_28_sva,
      regs_24_sva, regs_29_sva, regs_25_sva, {(MAC_and_43_nl) , (MAC_and_44_nl) ,
      (MAC_and_45_nl) , (MAC_and_46_nl) , (MAC_and_47_nl) , (MAC_and_48_nl) , (MAC_and_49_nl)});

  function automatic [0:0] MUX1HOT_s_1_15_2;
    input [0:0] input_14;
    input [0:0] input_13;
    input [0:0] input_12;
    input [0:0] input_11;
    input [0:0] input_10;
    input [0:0] input_9;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [14:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    result = result | ( input_9 & {1{sel[9]}});
    result = result | ( input_10 & {1{sel[10]}});
    result = result | ( input_11 & {1{sel[11]}});
    result = result | ( input_12 & {1{sel[12]}});
    result = result | ( input_13 & {1{sel[13]}});
    result = result | ( input_14 & {1{sel[14]}});
    MUX1HOT_s_1_15_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_6_2;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [5:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_9_2;
    input [0:0] input_8;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [8:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    result = result | ( input_8 & {1{sel[8]}});
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_4_2;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [3:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    MUX1HOT_v_16_4_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_7_2;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [6:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    result = result | ( input_5 & {16{sel[5]}});
    result = result | ( input_6 & {16{sel[6]}});
    MUX1HOT_v_16_7_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_3_2;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [2:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    MUX1HOT_v_30_3_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_5_2;
    input [29:0] input_4;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [4:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    result = result | ( input_3 & {30{sel[3]}});
    result = result | ( input_4 & {30{sel[4]}});
    MUX1HOT_v_30_5_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_6_2;
    input [29:0] input_5;
    input [29:0] input_4;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [5:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    result = result | ( input_3 & {30{sel[3]}});
    result = result | ( input_4 & {30{sel[4]}});
    result = result | ( input_5 & {30{sel[5]}});
    MUX1HOT_v_30_6_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_u2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_6 =  {1'b0, vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, coeffs_rsc_radr, coeffs_rsc_q, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz,
      out1_rsc_dat, out1_rsc_triosy_lz
);
  input clk;
  input rst;
  output [4:0] coeffs_rsc_radr;
  input [15:0] coeffs_rsc_q;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;


  // Interconnect Declarations
  wire [4:0] coeffs_rsci_radr_d;
  wire [15:0] coeffs_rsci_q_d;
  wire coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen coeffs_rsci (
      .q(coeffs_rsc_q),
      .radr(coeffs_rsc_radr),
      .radr_d(coeffs_rsci_radr_d),
      .q_d(coeffs_rsci_q_d),
      .rport_r_ram_ir_internal_RMASK_B_d(coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d)
    );
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .coeffs_rsc_triosy_lz(coeffs_rsc_triosy_lz),
      .in1_rsc_dat(in1_rsc_dat),
      .in1_rsc_triosy_lz(in1_rsc_triosy_lz),
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_triosy_lz(out1_rsc_triosy_lz),
      .coeffs_rsci_radr_d(coeffs_rsci_radr_d),
      .coeffs_rsci_q_d(coeffs_rsci_q_d),
      .coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d(coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d)
    );
endmodule



