
//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.3d/815731 Production Release
//  HLS Date:       Wed Apr 24 14:54:19 PDT 2019
// 
//  Generated by:   695r48@cparch23.ecn.purdue.edu
//  Generated date: Tue Nov  9 15:17:43 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen
// ------------------------------------------------------------------


module fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen (
  q, radr, radr_d, q_d, rport_r_ram_ir_internal_RMASK_B_d
);
  input [15:0] q;
  output [4:0] radr;
  input [4:0] radr_d;
  output [15:0] q_d;
  input rport_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_core_core_fsm (
  clk, rst, fsm_output, MAC_C_5_tr0
);
  input clk;
  input rst;
  output [18:0] fsm_output;
  reg [18:0] fsm_output;
  input MAC_C_5_tr0;


  // FSM State Type Declaration for fir_core_core_fsm_1
  parameter
    main_C_0 = 5'd0,
    MAC_C_0 = 5'd1,
    MAC_C_1 = 5'd2,
    MAC_C_2 = 5'd3,
    MAC_C_3 = 5'd4,
    MAC_C_4 = 5'd5,
    MAC_C_5 = 5'd6,
    MAC_C_6 = 5'd7,
    MAC_C_7 = 5'd8,
    MAC_C_8 = 5'd9,
    MAC_C_9 = 5'd10,
    MAC_C_10 = 5'd11,
    MAC_C_11 = 5'd12,
    MAC_C_12 = 5'd13,
    MAC_C_13 = 5'd14,
    MAC_C_14 = 5'd15,
    MAC_C_15 = 5'd16,
    MAC_C_16 = 5'd17,
    main_C_1 = 5'd18;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_core_core_fsm_1
    case (state_var)
      MAC_C_0 : begin
        fsm_output = 19'b0000000000000000010;
        state_var_NS = MAC_C_1;
      end
      MAC_C_1 : begin
        fsm_output = 19'b0000000000000000100;
        state_var_NS = MAC_C_2;
      end
      MAC_C_2 : begin
        fsm_output = 19'b0000000000000001000;
        state_var_NS = MAC_C_3;
      end
      MAC_C_3 : begin
        fsm_output = 19'b0000000000000010000;
        state_var_NS = MAC_C_4;
      end
      MAC_C_4 : begin
        fsm_output = 19'b0000000000000100000;
        state_var_NS = MAC_C_5;
      end
      MAC_C_5 : begin
        fsm_output = 19'b0000000000001000000;
        if ( MAC_C_5_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = MAC_C_6;
        end
      end
      MAC_C_6 : begin
        fsm_output = 19'b0000000000010000000;
        state_var_NS = MAC_C_7;
      end
      MAC_C_7 : begin
        fsm_output = 19'b0000000000100000000;
        state_var_NS = MAC_C_8;
      end
      MAC_C_8 : begin
        fsm_output = 19'b0000000001000000000;
        state_var_NS = MAC_C_9;
      end
      MAC_C_9 : begin
        fsm_output = 19'b0000000010000000000;
        state_var_NS = MAC_C_10;
      end
      MAC_C_10 : begin
        fsm_output = 19'b0000000100000000000;
        state_var_NS = MAC_C_11;
      end
      MAC_C_11 : begin
        fsm_output = 19'b0000001000000000000;
        state_var_NS = MAC_C_12;
      end
      MAC_C_12 : begin
        fsm_output = 19'b0000010000000000000;
        state_var_NS = MAC_C_13;
      end
      MAC_C_13 : begin
        fsm_output = 19'b0000100000000000000;
        state_var_NS = MAC_C_14;
      end
      MAC_C_14 : begin
        fsm_output = 19'b0001000000000000000;
        state_var_NS = MAC_C_15;
      end
      MAC_C_15 : begin
        fsm_output = 19'b0010000000000000000;
        state_var_NS = MAC_C_16;
      end
      MAC_C_16 : begin
        fsm_output = 19'b0100000000000000000;
        state_var_NS = MAC_C_0;
      end
      main_C_1 : begin
        fsm_output = 19'b1000000000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 19'b0000000000000000001;
        state_var_NS = MAC_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz, out1_rsc_dat, out1_rsc_triosy_lz,
      coeffs_rsci_radr_d, coeffs_rsci_q_d, coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d
);
  input clk;
  input rst;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;
  output [4:0] coeffs_rsci_radr_d;
  input [15:0] coeffs_rsci_q_d;
  output coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire [15:0] in1_rsci_idat;
  reg [15:0] out1_rsci_idat;
  wire [18:0] fsm_output;
  wire [4:0] MAC_acc_6_tmp;
  wire [5:0] nl_MAC_acc_6_tmp;
  wire and_dcpl_21;
  wire and_dcpl_22;
  wire and_dcpl_33;
  wire or_dcpl_26;
  wire or_dcpl_30;
  wire or_dcpl_31;
  wire or_dcpl_38;
  wire or_tmp_163;
  wire or_tmp_172;
  reg reg_out1_rsc_triosy_obj_ld_cse;
  wire reg_out1_out1_and_cse;
  wire coeffs_or_cse;
  wire coeffs_or_9_cse;
  wire nor_11_cse;
  reg [3:0] MAC_slc_MAC_2_MAC_acc_psp_sva;
  reg [1:0] MAC_acc_4_psp_sva;
  wire [2:0] nl_MAC_acc_4_psp_sva;
  reg [2:0] MAC_acc_psp_sva;
  wire [29:0] z_out_1;
  wire signed [31:0] nl_z_out_1;
  wire [29:0] z_out_2;
  wire signed [31:0] nl_z_out_2;
  wire [29:0] z_out_3;
  wire signed [31:0] nl_z_out_3;
  wire [29:0] z_out_4;
  wire signed [31:0] nl_z_out_4;
  wire [3:0] z_out_6;
  wire [4:0] nl_z_out_6;
  reg [15:0] regs_15_sva;
  reg [15:0] regs_16_sva;
  reg [15:0] regs_14_sva;
  reg [15:0] regs_17_sva;
  reg [15:0] regs_13_sva;
  reg [15:0] regs_18_sva;
  reg [15:0] regs_12_sva;
  reg [15:0] regs_19_sva;
  reg [15:0] regs_11_sva;
  reg [15:0] regs_20_sva;
  reg [15:0] regs_10_sva;
  reg [15:0] regs_21_sva;
  reg [15:0] regs_9_sva;
  reg [15:0] regs_22_sva;
  reg [15:0] regs_8_sva;
  reg [15:0] regs_23_sva;
  reg [15:0] regs_7_sva;
  reg [15:0] regs_24_sva;
  reg [15:0] regs_6_sva;
  reg [15:0] regs_25_sva;
  reg [15:0] regs_5_sva;
  reg [15:0] regs_26_sva;
  reg [15:0] regs_4_sva;
  reg [15:0] regs_27_sva;
  reg [15:0] regs_3_sva;
  reg [15:0] regs_28_sva;
  reg [15:0] regs_2_sva;
  reg [15:0] regs_29_sva;
  reg [15:0] regs_1_sva;
  reg [15:0] regs_30_sva;
  reg [15:0] regs_0_sva;
  reg [29:0] acc_32_3_1_sva;
  reg [15:0] regs_30_sva_1;
  reg [15:0] regs_29_sva_1;
  reg [15:0] regs_28_sva_1;
  reg [15:0] regs_27_sva_1;
  reg [15:0] regs_26_sva_1;
  reg [15:0] regs_25_sva_1;
  reg [15:0] regs_24_sva_1;
  reg [15:0] regs_23_sva_1;
  reg [15:0] regs_22_sva_1;
  reg [15:0] regs_21_sva_1;
  reg [15:0] regs_20_sva_1;
  reg [15:0] regs_19_sva_1;
  reg [15:0] regs_18_sva_1;
  reg [15:0] regs_17_sva_1;
  reg [15:0] regs_16_sva_1;
  reg [15:0] regs_15_sva_1;
  reg [15:0] regs_14_sva_1;
  reg [15:0] regs_13_sva_1;
  reg [15:0] regs_12_sva_1;
  reg [15:0] regs_11_sva_1;
  reg [15:0] regs_10_sva_1;
  reg [15:0] regs_9_sva_1;
  reg [15:0] regs_8_sva_1;
  reg [15:0] regs_7_sva_1;
  reg [15:0] regs_6_sva_1;
  reg [15:0] regs_5_sva_1;
  reg [15:0] regs_4_sva_1;
  reg [15:0] regs_3_sva_1;
  reg [15:0] regs_2_sva_1;
  reg [15:0] regs_1_sva_1;
  reg [15:0] regs_0_sva_1;
  reg [15:0] MAC_3_MAC_mux_itm;
  reg [15:0] MAC_4_MAC_mux_itm;
  reg [15:0] MAC_1_MAC_mux_itm;
  reg [15:0] MAC_9_MAC_mux_itm;
  reg [15:0] MAC_10_MAC_mux_itm;
  reg [29:0] MAC_10_mul_itm;
  reg [15:0] MAC_11_MAC_mux_itm;
  reg [29:0] MAC_11_mul_itm;
  reg [15:0] MAC_12_MAC_mux_itm;
  reg [29:0] MAC_acc_11_itm;
  reg [15:0] MAC_13_MAC_mux_itm;
  reg [15:0] MAC_14_MAC_mux_itm;
  reg [15:0] MAC_5_MAC_mux_itm;
  reg [15:0] MAC_6_MAC_mux_itm;
  reg [15:0] MAC_7_MAC_mux_itm;
  reg [15:0] MAC_8_MAC_mux_itm;
  reg [29:0] MAC_acc_17_itm;
  wire [29:0] MAC_acc_9_mx0w2;
  wire [30:0] nl_MAC_acc_9_mx0w2;
  wire [29:0] acc_32_3_5_sva_1;
  wire [30:0] nl_acc_32_3_5_sva_1;
  wire [3:0] MAC_slc_MAC_2_MAC_acc_psp_sva_mx0w0;
  wire [4:0] nl_MAC_slc_MAC_2_MAC_acc_psp_sva_mx0w0;
  wire [2:0] MAC_acc_psp_sva_1;
  wire [3:0] nl_MAC_acc_psp_sva_1;
  wire [29:0] MAC_acc_8_itm_mx0w0;
  wire [30:0] nl_MAC_acc_8_itm_mx0w0;
  wire [29:0] MAC_acc_16_mx0w0;
  wire [30:0] nl_MAC_acc_16_mx0w0;
  wire or_232_tmp;
  wire or_228_tmp;
  wire or_227_tmp;
  wire or_226_tmp;
  wire or_225_tmp;
  wire and_458_tmp;
  wire and_452_tmp;
  wire MAC_and_31_rgt;
  wire MAC_and_32_rgt;
  wire MAC_and_33_rgt;
  wire MAC_and_34_rgt;
  wire MAC_and_27_rgt;
  wire MAC_and_28_rgt;
  wire MAC_and_29_rgt;
  wire MAC_and_30_rgt;
  reg [1:0] MAC_i_5_1_sva_rsp_0;
  reg [1:0] MAC_i_5_1_sva_rsp_2;
  reg MAC_acc_3_psp_sva_rsp_0;
  reg MAC_acc_3_psp_sva_rsp_2;
  reg MAC_acc_5_itm_3;
  reg [1:0] MAC_acc_5_itm_2_1;
  reg MAC_acc_5_itm_0;
  wire MAC_nor_1_cse;
  wire MAC_i_or_2_cse;
  wire MAC_nor_2_cse;
  wire MAC_nor_3_cse;
  wire MAC_nor_4_cse;
  wire MAC_nor_8_cse;
  wire MAC_nor_9_cse;

  wire[29:0] acc_mux1h_1_nl;
  wire[29:0] MAC_14_acc_1_nl;
  wire[30:0] nl_MAC_14_acc_1_nl;
  wire[0:0] acc_not_nl;
  wire[0:0] MAC_i_MAC_i_mux_1_nl;
  wire[1:0] MAC_i_MAC_i_or_nl;
  wire[0:0] MAC_i_or_nl;
  wire[0:0] MAC_i_MAC_i_mux_nl;
  wire[0:0] MAC_and_38_nl;
  wire[0:0] MAC_and_36_nl;
  wire[0:0] MAC_MAC_nor_7_nl;
  wire[0:0] MAC_and_22_nl;
  wire[0:0] MAC_and_23_nl;
  wire[0:0] MAC_and_24_nl;
  wire[0:0] MAC_and_25_nl;
  wire[0:0] MAC_and_26_nl;
  wire[0:0] MAC_MAC_nor_8_nl;
  wire[0:0] MAC_and_16_nl;
  wire[0:0] MAC_and_17_nl;
  wire[0:0] MAC_and_18_nl;
  wire[0:0] MAC_and_19_nl;
  wire[0:0] MAC_and_20_nl;
  wire[0:0] MAC_and_14_nl;
  wire[0:0] MAC_and_12_nl;
  wire[0:0] MAC_and_nl;
  wire[0:0] MAC_and_1_nl;
  wire[0:0] MAC_and_2_nl;
  wire[0:0] MAC_and_7_nl;
  wire[0:0] MAC_and_8_nl;
  wire[0:0] MAC_and_9_nl;
  wire[0:0] MAC_and_10_nl;
  wire[0:0] MAC_and_3_nl;
  wire[0:0] MAC_and_4_nl;
  wire[0:0] MAC_and_5_nl;
  wire[0:0] MAC_and_6_nl;
  wire[29:0] mul_nl;
  wire signed [31:0] nl_mul_nl;
  wire[15:0] MAC_mux_31_nl;
  wire[0:0] MAC_or_nl;
  wire[0:0] MAC_or_4_nl;
  wire[29:0] mul_5_nl;
  wire signed [31:0] nl_mul_5_nl;
  wire[15:0] MAC_mux_36_nl;
  wire[29:0] MAC_3_mul_nl;
  wire signed [31:0] nl_MAC_3_mul_nl;
  wire[29:0] MAC_acc_18_nl;
  wire[30:0] nl_MAC_acc_18_nl;
  wire[0:0] MAC_or_2_nl;
  wire[0:0] coeffs_mux1h_1_nl;
  wire[0:0] coeffs_or_7_nl;
  wire[0:0] coeffs_or_1_nl;
  wire[2:0] coeffs_mux1h_2_nl;
  wire[0:0] coeffs_or_2_nl;
  wire[0:0] coeffs_or_3_nl;
  wire[0:0] coeffs_or_4_nl;
  wire[0:0] coeffs_or_5_nl;
  wire[0:0] coeffs_coeffs_or_nl;
  wire[15:0] MAC_mux_32_nl;
  wire[0:0] or_265_nl;
  wire[15:0] MAC_mux_33_nl;
  wire[15:0] MAC_mux_34_nl;
  wire[15:0] MAC_mux_35_nl;
  wire[0:0] MAC_mux_37_nl;
  wire[2:0] MAC_mux_38_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_fir_core_core_fsm_inst_MAC_C_5_tr0;
  assign nl_fir_core_core_fsm_inst_MAC_C_5_tr0 = MAC_i_5_1_sva_rsp_0[1];
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd16)) in1_rsci (
      .dat(in1_rsc_dat),
      .idat(in1_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd16)) out1_rsci (
      .idat(out1_rsci_idat),
      .dat(out1_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) coeffs_rsc_triosy_obj (
      .ld(reg_out1_rsc_triosy_obj_ld_cse),
      .lz(coeffs_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) in1_rsc_triosy_obj (
      .ld(reg_out1_rsc_triosy_obj_ld_cse),
      .lz(in1_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) out1_rsc_triosy_obj (
      .ld(reg_out1_rsc_triosy_obj_ld_cse),
      .lz(out1_rsc_triosy_lz)
    );
  fir_core_core_fsm fir_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .MAC_C_5_tr0(nl_fir_core_core_fsm_inst_MAC_C_5_tr0[0:0])
    );
  assign reg_out1_out1_and_cse = (fsm_output[6]) & (MAC_i_5_1_sva_rsp_0[1]);
  assign nor_11_cse = ~((fsm_output[18]) | (fsm_output[0]));
  assign MAC_i_or_2_cse = nor_11_cse & (~ (fsm_output[2]));
  assign MAC_nor_1_cse = ~((MAC_acc_psp_sva_1[1:0]!=2'b00));
  assign MAC_and_31_rgt = ~((z_out_6[3]) | (z_out_6[0]) | and_458_tmp);
  assign MAC_and_32_rgt = (z_out_6[0]) & (~ (z_out_6[3])) & (~ and_458_tmp);
  assign MAC_and_33_rgt = (z_out_6[3]) & (~ (z_out_6[0])) & (~ and_458_tmp);
  assign MAC_and_34_rgt = (z_out_6[3]) & (z_out_6[0]) & (~ and_458_tmp);
  assign MAC_and_27_rgt = ~((z_out_6[3]) | (z_out_6[0]) | or_tmp_172);
  assign MAC_and_28_rgt = (z_out_6[0]) & (~ (z_out_6[3])) & (~ or_tmp_172);
  assign MAC_and_29_rgt = (z_out_6[3]) & (~ (z_out_6[0])) & (~ or_tmp_172);
  assign MAC_and_30_rgt = (z_out_6[3]) & (z_out_6[0]) & (~ or_tmp_172);
  assign MAC_nor_2_cse = ~((MAC_acc_6_tmp[3]) | (MAC_acc_6_tmp[1]));
  assign MAC_nor_3_cse = ~((MAC_acc_6_tmp[3]) | (MAC_acc_6_tmp[0]));
  assign MAC_nor_4_cse = ~((MAC_acc_6_tmp[1:0]!=2'b00));
  assign MAC_nor_8_cse = ~(MAC_acc_3_psp_sva_rsp_0 | (MAC_acc_4_psp_sva[1]));
  assign MAC_nor_9_cse = ~(MAC_acc_3_psp_sva_rsp_0 | (MAC_acc_4_psp_sva[0]));
  assign nl_MAC_acc_9_mx0w2 = MAC_acc_8_itm_mx0w0 + acc_32_3_1_sva;
  assign MAC_acc_9_mx0w2 = nl_MAC_acc_9_mx0w2[29:0];
  assign nl_acc_32_3_5_sva_1 = MAC_acc_9_mx0w2 + MAC_acc_11_itm;
  assign acc_32_3_5_sva_1 = nl_acc_32_3_5_sva_1[29:0];
  assign nl_MAC_acc_6_tmp = conv_u2s_4_5(MAC_slc_MAC_2_MAC_acc_psp_sva_mx0w0) + 5'b00001;
  assign MAC_acc_6_tmp = nl_MAC_acc_6_tmp[4:0];
  assign nl_MAC_slc_MAC_2_MAC_acc_psp_sva_mx0w0 = ({MAC_acc_5_itm_3 , MAC_acc_5_itm_2_1
      , MAC_acc_5_itm_0}) + 4'b0001;
  assign MAC_slc_MAC_2_MAC_acc_psp_sva_mx0w0 = nl_MAC_slc_MAC_2_MAC_acc_psp_sva_mx0w0[3:0];
  assign nl_MAC_acc_psp_sva_1 = conv_u2u_2_3({1'b1 , (~ (MAC_acc_6_tmp[0]))}) + 3'b001;
  assign MAC_acc_psp_sva_1 = nl_MAC_acc_psp_sva_1[2:0];
  assign nl_MAC_acc_8_itm_mx0w0 = MAC_11_mul_itm + MAC_10_mul_itm;
  assign MAC_acc_8_itm_mx0w0 = nl_MAC_acc_8_itm_mx0w0[29:0];
  assign nl_MAC_acc_16_mx0w0 = MAC_acc_8_itm_mx0w0 + MAC_acc_11_itm;
  assign MAC_acc_16_mx0w0 = nl_MAC_acc_16_mx0w0[29:0];
  assign and_dcpl_21 = ~((fsm_output[17:16]!=2'b00));
  assign and_dcpl_22 = and_dcpl_21 & (~ (fsm_output[15]));
  assign and_dcpl_33 = ~((fsm_output[1]) | (fsm_output[14]));
  assign or_dcpl_26 = (fsm_output[8]) | (fsm_output[6]);
  assign or_dcpl_30 = (fsm_output[5:4]!=2'b00);
  assign or_dcpl_31 = or_dcpl_30 | (fsm_output[3]) | (fsm_output[7]);
  assign or_dcpl_38 = or_dcpl_30 | (fsm_output[3]);
  assign or_tmp_163 = ~((~ and_dcpl_21) | (fsm_output[15]) | (fsm_output[18]) | (fsm_output[0])
      | (fsm_output[1]) | (fsm_output[14]));
  assign or_tmp_172 = and_dcpl_22 & (~ (fsm_output[13])) & (~ (fsm_output[18])) &
      (~ (fsm_output[0])) & (~ (fsm_output[12])) & and_dcpl_33;
  assign coeffs_or_cse = (fsm_output[2:1]!=2'b00);
  assign coeffs_or_9_cse = (fsm_output[4:3]!=2'b00);
  assign coeffs_or_7_nl = (fsm_output[5]) | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[13])
      | (fsm_output[14]);
  assign coeffs_or_1_nl = (fsm_output[12:9]!=4'b0000);
  assign coeffs_mux1h_1_nl = MUX1HOT_s_1_5_2(MAC_acc_5_itm_3, (MAC_slc_MAC_2_MAC_acc_psp_sva[3]),
      (MAC_i_5_1_sva_rsp_0[0]), (MAC_i_5_1_sva_rsp_0[0]), MAC_acc_3_psp_sva_rsp_0,
      {coeffs_or_cse , coeffs_or_9_cse , (coeffs_or_7_nl) , (fsm_output[6]) , (coeffs_or_1_nl)});
  assign coeffs_or_2_nl = (fsm_output[8:7]!=2'b00);
  assign coeffs_or_3_nl = (fsm_output[10:9]!=2'b00);
  assign coeffs_or_4_nl = (fsm_output[12:11]!=2'b00);
  assign coeffs_or_5_nl = (fsm_output[14:13]!=2'b00);
  assign coeffs_mux1h_2_nl = MUX1HOT_v_3_8_2(({MAC_acc_5_itm_2_1 , MAC_acc_5_itm_0}),
      (MAC_slc_MAC_2_MAC_acc_psp_sva[2:0]), ({2'b01 , (~ (MAC_i_5_1_sva_rsp_2[0]))}),
      ({2'b01 , (~ (MAC_i_5_1_sva_rsp_2[0]))}), ({1'b0 , MAC_i_5_1_sva_rsp_2}), ({1'b1
      , MAC_acc_4_psp_sva}), ({2'b10 , MAC_acc_3_psp_sva_rsp_2}), MAC_acc_psp_sva,
      {coeffs_or_cse , coeffs_or_9_cse , (fsm_output[5]) , (fsm_output[6]) , (coeffs_or_2_nl)
      , (coeffs_or_3_nl) , (coeffs_or_4_nl) , (coeffs_or_5_nl)});
  assign coeffs_coeffs_or_nl = (fsm_output[1]) | (fsm_output[3]) | (fsm_output[5])
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[11]) | (fsm_output[13]);
  assign coeffs_rsci_radr_d = {(coeffs_mux1h_1_nl) , (coeffs_mux1h_2_nl) , (coeffs_coeffs_or_nl)};
  assign coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d = (and_dcpl_22 & nor_11_cse
      & (~ (fsm_output[6]))) | ((~ (MAC_i_5_1_sva_rsp_0[1])) & (fsm_output[6]));
  assign and_452_tmp = and_dcpl_22 & nor_11_cse & (~ (fsm_output[1]));
  assign and_458_tmp = and_dcpl_21 & (~ (fsm_output[15])) & (~ (fsm_output[13]))
      & nor_11_cse & and_dcpl_33;
  assign or_225_tmp = or_dcpl_31 | (fsm_output[2]) | (fsm_output[8]) | (fsm_output[6]);
  assign or_226_tmp = or_dcpl_38 | (fsm_output[7]) | (fsm_output[2]) | (fsm_output[6]);
  assign or_227_tmp = or_dcpl_38 | (fsm_output[2]) | (fsm_output[6]);
  assign or_228_tmp = or_dcpl_30 | (fsm_output[3:2]!=2'b00);
  assign or_232_tmp = or_dcpl_31 | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[6]);
  always @(posedge clk) begin
    if ( rst ) begin
      acc_32_3_1_sva <= 30'b000000000000000000000000000000;
    end
    else if ( (fsm_output[17]) | (fsm_output[0]) | (fsm_output[12]) | (fsm_output[6])
        ) begin
      acc_32_3_1_sva <= MUX_v_30_2_2(30'b000000000000000000000000000000, (acc_mux1h_1_nl),
          (acc_not_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out1_rsci_idat <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
      regs_14_sva <= 16'b0000000000000000;
      regs_28_sva <= 16'b0000000000000000;
      regs_13_sva <= 16'b0000000000000000;
      regs_27_sva <= 16'b0000000000000000;
      regs_2_sva <= 16'b0000000000000000;
      regs_16_sva <= 16'b0000000000000000;
      regs_30_sva <= 16'b0000000000000000;
      regs_1_sva <= 16'b0000000000000000;
      regs_15_sva <= 16'b0000000000000000;
      regs_29_sva <= 16'b0000000000000000;
      regs_10_sva <= 16'b0000000000000000;
      regs_12_sva <= 16'b0000000000000000;
      regs_26_sva <= 16'b0000000000000000;
      regs_9_sva <= 16'b0000000000000000;
      regs_11_sva <= 16'b0000000000000000;
      regs_25_sva <= 16'b0000000000000000;
      regs_6_sva <= 16'b0000000000000000;
      regs_20_sva <= 16'b0000000000000000;
      regs_5_sva <= 16'b0000000000000000;
      regs_19_sva <= 16'b0000000000000000;
      regs_4_sva <= 16'b0000000000000000;
      regs_18_sva <= 16'b0000000000000000;
      regs_3_sva <= 16'b0000000000000000;
      regs_17_sva <= 16'b0000000000000000;
      regs_8_sva <= 16'b0000000000000000;
      regs_24_sva <= 16'b0000000000000000;
      regs_7_sva <= 16'b0000000000000000;
      regs_23_sva <= 16'b0000000000000000;
      regs_22_sva <= 16'b0000000000000000;
      regs_21_sva <= 16'b0000000000000000;
    end
    else if ( reg_out1_out1_and_cse ) begin
      out1_rsci_idat <= acc_32_3_5_sva_1[29:14];
      regs_0_sva <= regs_0_sva_1;
      regs_14_sva <= regs_14_sva_1;
      regs_28_sva <= regs_28_sva_1;
      regs_13_sva <= regs_13_sva_1;
      regs_27_sva <= regs_27_sva_1;
      regs_2_sva <= regs_2_sva_1;
      regs_16_sva <= regs_16_sva_1;
      regs_30_sva <= regs_30_sva_1;
      regs_1_sva <= regs_1_sva_1;
      regs_15_sva <= regs_15_sva_1;
      regs_29_sva <= regs_29_sva_1;
      regs_10_sva <= regs_10_sva_1;
      regs_12_sva <= regs_12_sva_1;
      regs_26_sva <= regs_26_sva_1;
      regs_9_sva <= regs_9_sva_1;
      regs_11_sva <= regs_11_sva_1;
      regs_25_sva <= regs_25_sva_1;
      regs_6_sva <= regs_6_sva_1;
      regs_20_sva <= regs_20_sva_1;
      regs_5_sva <= regs_5_sva_1;
      regs_19_sva <= regs_19_sva_1;
      regs_4_sva <= regs_4_sva_1;
      regs_18_sva <= regs_18_sva_1;
      regs_3_sva <= regs_3_sva_1;
      regs_17_sva <= regs_17_sva_1;
      regs_8_sva <= regs_8_sva_1;
      regs_24_sva <= regs_24_sva_1;
      regs_7_sva <= regs_7_sva_1;
      regs_23_sva <= regs_23_sva_1;
      regs_22_sva <= regs_22_sva_1;
      regs_21_sva <= regs_21_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_0_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_0_sva_1 <= in1_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_out1_rsc_triosy_obj_ld_cse <= 1'b0;
      MAC_acc_5_itm_3 <= 1'b0;
      MAC_acc_5_itm_2_1 <= 2'b00;
      MAC_acc_5_itm_0 <= 1'b0;
      MAC_11_mul_itm <= 30'b000000000000000000000000000000;
    end
    else begin
      reg_out1_rsc_triosy_obj_ld_cse <= reg_out1_out1_and_cse;
      MAC_acc_5_itm_3 <= (MAC_i_MAC_i_mux_1_nl) & nor_11_cse;
      MAC_acc_5_itm_2_1 <= MUX_v_2_2_2(2'b00, (MAC_i_MAC_i_or_nl), nor_11_cse);
      MAC_acc_5_itm_0 <= (MAC_i_MAC_i_mux_nl) & nor_11_cse;
      MAC_11_mul_itm <= MUX1HOT_v_30_7_2((mul_5_nl), (MAC_3_mul_nl), z_out_4, z_out_1,
          z_out_3, z_out_2, (MAC_acc_18_nl), {(MAC_or_2_nl) , (fsm_output[5]) , (fsm_output[9])
          , (fsm_output[11]) , (fsm_output[13]) , (fsm_output[15]) , (fsm_output[16])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_30_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_30_sva_1 <= regs_29_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_29_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_29_sva_1 <= regs_28_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_28_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_28_sva_1 <= regs_27_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_27_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_27_sva_1 <= regs_26_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_26_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_26_sva_1 <= regs_25_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_25_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_25_sva_1 <= regs_24_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_24_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_24_sva_1 <= regs_23_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_23_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_23_sva_1 <= regs_22_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_22_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_22_sva_1 <= regs_21_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_21_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_21_sva_1 <= regs_20_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_20_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_20_sva_1 <= regs_19_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_19_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_19_sva_1 <= regs_18_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_18_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_18_sva_1 <= regs_17_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_17_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_17_sva_1 <= regs_16_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_16_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_16_sva_1 <= regs_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_15_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_15_sva_1 <= regs_14_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_14_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_14_sva_1 <= regs_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_13_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_13_sva_1 <= regs_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_12_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_12_sva_1 <= regs_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_11_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_11_sva_1 <= regs_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_10_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_10_sva_1 <= regs_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_9_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_9_sva_1 <= regs_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_8_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_8_sva_1 <= regs_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_7_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_7_sva_1 <= regs_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_6_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_6_sva_1 <= regs_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_5_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_5_sva_1 <= regs_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_4_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_4_sva_1 <= regs_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_3_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_3_sva_1 <= regs_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_2_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_2_sva_1 <= regs_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      regs_1_sva_1 <= 16'b0000000000000000;
    end
    else if ( ~ nor_11_cse ) begin
      regs_1_sva_1 <= regs_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_3_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( fsm_output[1] ) begin
      MAC_3_MAC_mux_itm <= MUX_v_16_16_2x0x2x3x4x5x6x7x9x10x11x12x13x14(regs_1_sva,
          regs_15_sva, regs_29_sva, MAC_slc_MAC_2_MAC_acc_psp_sva_mx0w0);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_4_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( fsm_output[1] ) begin
      MAC_4_MAC_mux_itm <= MUX_v_16_16_2x0x2x3x4x5x6x7x9x10x11x12x13x14(regs_2_sva,
          regs_16_sva, regs_30_sva, MAC_slc_MAC_2_MAC_acc_psp_sva_mx0w0);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_slc_MAC_2_MAC_acc_psp_sva <= 4'b0000;
    end
    else if ( fsm_output[1] ) begin
      MAC_slc_MAC_2_MAC_acc_psp_sva <= MAC_slc_MAC_2_MAC_acc_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( fsm_output[1] ) begin
      MAC_1_MAC_mux_itm <= MUX_v_16_15_2x1x2x3x4x5x6x8x9x10x11x12x13(regs_0_sva_1,
          regs_13_sva, regs_27_sva, {MAC_acc_5_itm_3 , MAC_acc_5_itm_2_1 , MAC_acc_5_itm_0});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_9_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ and_452_tmp ) begin
      MAC_9_MAC_mux_itm <= MUX_v_16_2_2(regs_21_sva, regs_7_sva, MAC_and_38_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_10_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_tmp_163 ) begin
      MAC_10_MAC_mux_itm <= MUX_v_16_2_2(regs_22_sva, regs_8_sva, MAC_and_36_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_psp_sva <= 3'b000;
    end
    else if ( ~ or_tmp_163 ) begin
      MAC_acc_psp_sva <= MAC_acc_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_11_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( MAC_and_31_rgt | MAC_and_32_rgt | MAC_and_33_rgt | MAC_and_34_rgt )
        begin
      MAC_11_MAC_mux_itm <= MUX1HOT_v_16_4_2(regs_7_sva, regs_9_sva, regs_23_sva,
          regs_25_sva, {MAC_and_31_rgt , MAC_and_32_rgt , MAC_and_33_rgt , MAC_and_34_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_12_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( MAC_and_27_rgt | MAC_and_28_rgt | MAC_and_29_rgt | MAC_and_30_rgt )
        begin
      MAC_12_MAC_mux_itm <= MUX1HOT_v_16_4_2(regs_8_sva, regs_10_sva, regs_24_sva,
          regs_26_sva, {MAC_and_27_rgt , MAC_and_28_rgt , MAC_and_29_rgt , MAC_and_30_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_4_psp_sva <= 2'b00;
    end
    else if ( ~(or_dcpl_31 | (fsm_output[9]) | (fsm_output[2]) | or_dcpl_26) ) begin
      MAC_acc_4_psp_sva <= nl_MAC_acc_4_psp_sva[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_5_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_225_tmp ) begin
      MAC_5_MAC_mux_itm <= MUX1HOT_v_16_6_2(regs_0_sva_1, regs_1_sva, regs_3_sva,
          regs_15_sva, regs_17_sva, regs_19_sva, {(MAC_MAC_nor_7_nl) , (MAC_and_22_nl)
          , (MAC_and_23_nl) , (MAC_and_24_nl) , (MAC_and_25_nl) , (MAC_and_26_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_6_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_226_tmp ) begin
      MAC_6_MAC_mux_itm <= MUX1HOT_v_16_6_2(regs_0_sva, regs_2_sva, regs_4_sva, regs_16_sva,
          regs_18_sva, regs_20_sva, {(MAC_MAC_nor_8_nl) , (MAC_and_16_nl) , (MAC_and_17_nl)
          , (MAC_and_18_nl) , (MAC_and_19_nl) , (MAC_and_20_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_7_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_227_tmp ) begin
      MAC_7_MAC_mux_itm <= MUX_v_16_2_2(regs_5_sva, regs_19_sva, MAC_and_14_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_228_tmp ) begin
      MAC_8_MAC_mux_itm <= MUX_v_16_2_2(regs_6_sva, regs_20_sva, MAC_and_12_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_13_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~(or_dcpl_31 | (fsm_output[10:9]!=2'b00) | or_dcpl_26) ) begin
      MAC_13_MAC_mux_itm <= MUX1HOT_v_16_7_2(regs_0_sva, regs_14_sva, regs_28_sva,
          regs_9_sva, regs_11_sva, regs_25_sva, regs_27_sva, {(MAC_and_nl) , (MAC_and_1_nl)
          , (MAC_and_2_nl) , (MAC_and_7_nl) , (MAC_and_8_nl) , (MAC_and_9_nl) , (MAC_and_10_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_MAC_mux_itm <= 16'b0000000000000000;
    end
    else if ( ~ or_232_tmp ) begin
      MAC_14_MAC_mux_itm <= MUX1HOT_v_16_4_2(regs_10_sva, regs_12_sva, regs_26_sva,
          regs_28_sva, {(MAC_and_3_nl) , (MAC_and_4_nl) , (MAC_and_5_nl) , (MAC_and_6_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_10_mul_itm <= 30'b000000000000000000000000000000;
    end
    else if ( (fsm_output[4]) | (fsm_output[12]) | (fsm_output[10]) | (fsm_output[2])
        | (fsm_output[14]) | (fsm_output[8]) | (fsm_output[6]) ) begin
      MAC_10_mul_itm <= MUX1HOT_v_30_5_2(z_out_1, (mul_nl), z_out_2, z_out_3, z_out_4,
          {(MAC_or_nl) , (MAC_or_4_nl) , (fsm_output[10]) , (fsm_output[12]) , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_11_itm <= 30'b000000000000000000000000000000;
    end
    else if ( (fsm_output[4]) | (fsm_output[14]) | (fsm_output[8]) ) begin
      MAC_acc_11_itm <= MAC_acc_8_itm_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_17_itm <= 30'b000000000000000000000000000000;
    end
    else if ( fsm_output[10] ) begin
      MAC_acc_17_itm <= MAC_acc_16_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_i_5_1_sva_rsp_0 <= 2'b00;
    end
    else if ( ~ or_tmp_163 ) begin
      MAC_i_5_1_sva_rsp_0 <= MAC_acc_6_tmp[4:3];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_i_5_1_sva_rsp_2 <= 2'b00;
    end
    else if ( ~ or_tmp_163 ) begin
      MAC_i_5_1_sva_rsp_2 <= MAC_acc_6_tmp[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_3_psp_sva_rsp_0 <= 1'b0;
    end
    else if ( ~ or_tmp_172 ) begin
      MAC_acc_3_psp_sva_rsp_0 <= z_out_6[3];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_acc_3_psp_sva_rsp_2 <= 1'b0;
    end
    else if ( ~ or_tmp_172 ) begin
      MAC_acc_3_psp_sva_rsp_2 <= z_out_6[0];
    end
  end
  assign nl_MAC_14_acc_1_nl = MAC_11_mul_itm + MAC_acc_17_itm;
  assign MAC_14_acc_1_nl = nl_MAC_14_acc_1_nl[29:0];
  assign acc_mux1h_1_nl = MUX1HOT_v_30_3_2(acc_32_3_5_sva_1, MAC_acc_9_mx0w2, (MAC_14_acc_1_nl),
      {(fsm_output[6]) , (fsm_output[12]) , (fsm_output[17])});
  assign acc_not_nl = ~ (fsm_output[0]);
  assign MAC_i_MAC_i_mux_1_nl = MUX_s_1_2_2((z_out_6[3]), MAC_acc_5_itm_3, MAC_i_or_2_cse);
  assign MAC_i_or_nl = (fsm_output[2]) | (fsm_output[6]);
  assign MAC_i_MAC_i_or_nl = MUX_v_2_2_2(MAC_acc_5_itm_2_1, 2'b11, (MAC_i_or_nl));
  assign MAC_i_MAC_i_mux_nl = MUX_s_1_2_2((z_out_6[0]), MAC_acc_5_itm_0, MAC_i_or_2_cse);
  assign MAC_mux_36_nl = MUX_v_16_2_2(MAC_1_MAC_mux_itm, MAC_7_MAC_mux_itm, fsm_output[7]);
  assign nl_mul_5_nl = $signed((MAC_mux_36_nl)) * $signed((coeffs_rsci_q_d));
  assign mul_5_nl = nl_mul_5_nl[29:0];
  assign nl_MAC_3_mul_nl = $signed(MAC_3_MAC_mux_itm) * $signed((coeffs_rsci_q_d));
  assign MAC_3_mul_nl = nl_MAC_3_mul_nl[29:0];
  assign nl_MAC_acc_18_nl = MAC_acc_16_mx0w0 + acc_32_3_1_sva;
  assign MAC_acc_18_nl = nl_MAC_acc_18_nl[29:0];
  assign MAC_or_2_nl = (fsm_output[3]) | (fsm_output[7]);
  assign MAC_and_38_nl = (MAC_acc_psp_sva_1[2]) & MAC_nor_1_cse & (~ and_452_tmp);
  assign MAC_and_36_nl = (MAC_acc_psp_sva_1[2]) & MAC_nor_1_cse & (~ or_tmp_163);
  assign nl_MAC_acc_4_psp_sva  = conv_u2u_1_2(z_out_6[0]) + 2'b01;
  assign MAC_MAC_nor_7_nl = ~((MAC_acc_6_tmp[3]) | (MAC_acc_6_tmp[1]) | (MAC_acc_6_tmp[0])
      | or_225_tmp);
  assign MAC_and_22_nl = (MAC_acc_6_tmp[0]) & MAC_nor_2_cse & (~ or_225_tmp);
  assign MAC_and_23_nl = (MAC_acc_6_tmp[1]) & MAC_nor_3_cse & (~ or_225_tmp);
  assign MAC_and_24_nl = (MAC_acc_6_tmp[3]) & MAC_nor_4_cse & (~ or_225_tmp);
  assign MAC_and_25_nl = (MAC_acc_6_tmp[3]) & (MAC_acc_6_tmp[0]) & (~ (MAC_acc_6_tmp[1]))
      & (~ or_225_tmp);
  assign MAC_and_26_nl = (MAC_acc_6_tmp[3]) & (MAC_acc_6_tmp[1]) & (~ (MAC_acc_6_tmp[0]))
      & (~ or_225_tmp);
  assign MAC_MAC_nor_8_nl = ~((MAC_acc_6_tmp[3]) | (MAC_acc_6_tmp[1]) | (MAC_acc_6_tmp[0])
      | or_226_tmp);
  assign MAC_and_16_nl = (MAC_acc_6_tmp[0]) & MAC_nor_2_cse & (~ or_226_tmp);
  assign MAC_and_17_nl = (MAC_acc_6_tmp[1]) & MAC_nor_3_cse & (~ or_226_tmp);
  assign MAC_and_18_nl = (MAC_acc_6_tmp[3]) & MAC_nor_4_cse & (~ or_226_tmp);
  assign MAC_and_19_nl = (MAC_acc_6_tmp[3]) & (MAC_acc_6_tmp[0]) & (~ (MAC_acc_6_tmp[1]))
      & (~ or_226_tmp);
  assign MAC_and_20_nl = (MAC_acc_6_tmp[3]) & (MAC_acc_6_tmp[1]) & (~ (MAC_acc_6_tmp[0]))
      & (~ or_226_tmp);
  assign MAC_and_14_nl = (MAC_acc_6_tmp[0]) & (~ or_227_tmp);
  assign MAC_and_12_nl = (MAC_acc_6_tmp[0]) & (~ or_228_tmp);
  assign MAC_and_nl = (~(MAC_acc_5_itm_3 | (MAC_acc_5_itm_2_1!=2'b00) | MAC_acc_5_itm_0))
      & (fsm_output[1]);
  assign MAC_and_1_nl = (MAC_acc_5_itm_2_1==2'b11) & MAC_acc_5_itm_0 & (~ MAC_acc_5_itm_3)
      & (fsm_output[1]);
  assign MAC_and_2_nl = MAC_acc_5_itm_3 & (MAC_acc_5_itm_2_1==2'b11) & (~ MAC_acc_5_itm_0)
      & (fsm_output[1]);
  assign MAC_and_7_nl = (MAC_acc_4_psp_sva[0]) & MAC_nor_8_cse & (fsm_output[2]);
  assign MAC_and_8_nl = (MAC_acc_4_psp_sva[1]) & MAC_nor_9_cse & (fsm_output[2]);
  assign MAC_and_9_nl = MAC_acc_3_psp_sva_rsp_0 & (MAC_acc_4_psp_sva==2'b01) & (fsm_output[2]);
  assign MAC_and_10_nl = MAC_acc_3_psp_sva_rsp_0 & (MAC_acc_4_psp_sva==2'b10) & (fsm_output[2]);
  assign MAC_and_3_nl = (MAC_acc_4_psp_sva[0]) & MAC_nor_8_cse & (~ or_232_tmp);
  assign MAC_and_4_nl = (MAC_acc_4_psp_sva[1]) & MAC_nor_9_cse & (~ or_232_tmp);
  assign MAC_and_5_nl = MAC_acc_3_psp_sva_rsp_0 & (MAC_acc_4_psp_sva==2'b01) & (~
      or_232_tmp);
  assign MAC_and_6_nl = MAC_acc_3_psp_sva_rsp_0 & (MAC_acc_4_psp_sva==2'b10) & (~
      or_232_tmp);
  assign MAC_mux_31_nl = MUX_v_16_2_2(MAC_4_MAC_mux_itm, MAC_8_MAC_mux_itm, fsm_output[6]);
  assign nl_mul_nl = $signed((MAC_mux_31_nl)) * $signed((coeffs_rsci_q_d));
  assign mul_nl = nl_mul_nl[29:0];
  assign MAC_or_nl = (fsm_output[2]) | (fsm_output[8]);
  assign MAC_or_4_nl = (fsm_output[4]) | (fsm_output[6]);
  assign or_265_nl = (fsm_output[11]) | (fsm_output[2]);
  assign MAC_mux_32_nl = MUX_v_16_2_2(MAC_6_MAC_mux_itm, MAC_13_MAC_mux_itm, or_265_nl);
  assign nl_z_out_1 = $signed((MAC_mux_32_nl)) * $signed((coeffs_rsci_q_d));
  assign z_out_1 = nl_z_out_1[29:0];
  assign MAC_mux_33_nl = MUX_v_16_2_2(MAC_14_MAC_mux_itm, MAC_9_MAC_mux_itm, fsm_output[15]);
  assign nl_z_out_2 = $signed((MAC_mux_33_nl)) * $signed((coeffs_rsci_q_d));
  assign z_out_2 = nl_z_out_2[29:0];
  assign MAC_mux_34_nl = MUX_v_16_2_2(MAC_12_MAC_mux_itm, MAC_11_MAC_mux_itm, fsm_output[13]);
  assign nl_z_out_3 = $signed((MAC_mux_34_nl)) * $signed((coeffs_rsci_q_d));
  assign z_out_3 = nl_z_out_3[29:0];
  assign MAC_mux_35_nl = MUX_v_16_2_2(MAC_10_MAC_mux_itm, MAC_5_MAC_mux_itm, fsm_output[9]);
  assign nl_z_out_4 = $signed((MAC_mux_35_nl)) * $signed((coeffs_rsci_q_d));
  assign z_out_4 = nl_z_out_4[29:0];
  assign MAC_mux_37_nl = MUX_s_1_2_2(MAC_acc_3_psp_sva_rsp_0, (MAC_acc_6_tmp[3]),
      fsm_output[1]);
  assign MAC_mux_38_nl = MUX_v_3_2_2(({1'b1 , MAC_acc_4_psp_sva}), MAC_acc_psp_sva_1,
      fsm_output[1]);
  assign nl_z_out_6 = ({(MAC_mux_37_nl) , (MAC_mux_38_nl)}) + 4'b0001;
  assign z_out_6 = nl_z_out_6[3:0];

  function automatic [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_4_2;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [3:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    MUX1HOT_v_16_4_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_6_2;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [5:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    result = result | ( input_5 & {16{sel[5]}});
    MUX1HOT_v_16_6_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_7_2;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [6:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    result = result | ( input_5 & {16{sel[5]}});
    result = result | ( input_6 & {16{sel[6]}});
    MUX1HOT_v_16_7_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_3_2;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [2:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    MUX1HOT_v_30_3_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_5_2;
    input [29:0] input_4;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [4:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    result = result | ( input_3 & {30{sel[3]}});
    result = result | ( input_4 & {30{sel[4]}});
    MUX1HOT_v_30_5_2 = result;
  end
  endfunction


  function automatic [29:0] MUX1HOT_v_30_7_2;
    input [29:0] input_6;
    input [29:0] input_5;
    input [29:0] input_4;
    input [29:0] input_3;
    input [29:0] input_2;
    input [29:0] input_1;
    input [29:0] input_0;
    input [6:0] sel;
    reg [29:0] result;
  begin
    result = input_0 & {30{sel[0]}};
    result = result | ( input_1 & {30{sel[1]}});
    result = result | ( input_2 & {30{sel[2]}});
    result = result | ( input_3 & {30{sel[3]}});
    result = result | ( input_4 & {30{sel[4]}});
    result = result | ( input_5 & {30{sel[5]}});
    result = result | ( input_6 & {30{sel[6]}});
    MUX1HOT_v_30_7_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_8_2;
    input [2:0] input_7;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [7:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    result = result | ( input_4 & {3{sel[4]}});
    result = result | ( input_5 & {3{sel[5]}});
    result = result | ( input_6 & {3{sel[6]}});
    result = result | ( input_7 & {3{sel[7]}});
    MUX1HOT_v_3_8_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_15_2x1x2x3x4x5x6x8x9x10x11x12x13;
    input [15:0] input_0;
    input [15:0] input_7;
    input [15:0] input_14;
    input [3:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0111 : begin
        result = input_7;
      end
      default : begin
        result = input_14;
      end
    endcase
    MUX_v_16_15_2x1x2x3x4x5x6x8x9x10x11x12x13 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_16_2x0x2x3x4x5x6x7x9x10x11x12x13x14;
    input [15:0] input_1;
    input [15:0] input_8;
    input [15:0] input_15;
    input [3:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      4'b0001 : begin
        result = input_1;
      end
      4'b1000 : begin
        result = input_8;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_16_16_2x0x2x3x4x5x6x7x9x10x11x12x13x14 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, coeffs_rsc_radr, coeffs_rsc_q, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz,
      out1_rsc_dat, out1_rsc_triosy_lz
);
  input clk;
  input rst;
  output [4:0] coeffs_rsc_radr;
  input [15:0] coeffs_rsc_q;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;


  // Interconnect Declarations
  wire [4:0] coeffs_rsci_radr_d;
  wire [15:0] coeffs_rsci_q_d;
  wire coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  fir_Altera_DIST_DIST_1R1W_RBW_rport_1_16_5_32_32_16_gen coeffs_rsci (
      .q(coeffs_rsc_q),
      .radr(coeffs_rsc_radr),
      .radr_d(coeffs_rsci_radr_d),
      .q_d(coeffs_rsci_q_d),
      .rport_r_ram_ir_internal_RMASK_B_d(coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d)
    );
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .coeffs_rsc_triosy_lz(coeffs_rsc_triosy_lz),
      .in1_rsc_dat(in1_rsc_dat),
      .in1_rsc_triosy_lz(in1_rsc_triosy_lz),
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_triosy_lz(out1_rsc_triosy_lz),
      .coeffs_rsci_radr_d(coeffs_rsci_radr_d),
      .coeffs_rsci_q_d(coeffs_rsci_q_d),
      .coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d(coeffs_rsci_rport_r_ram_ir_internal_RMASK_B_d)
    );
endmodule



