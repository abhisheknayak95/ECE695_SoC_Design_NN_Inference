
//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/mgc_in_wire_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_wire_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule


//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /package/eda/mg/Catapult_10.3d/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.3d/815731 Production Release
//  HLS Date:       Wed Apr 24 14:54:19 PDT 2019
// 
//  Generated by:   695r48@ecegrid-thin4.ecn.purdue.edu
//  Generated date: Wed Nov 10 16:27:37 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, coeffs_rsc_z, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz, out1_rsc_dat,
      out1_rsc_triosy_lz
);
  input clk;
  input rst;
  input [511:0] coeffs_rsc_z;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;


  // Interconnect Declarations
  wire [511:0] coeffs_rsci_d;
  wire [15:0] in1_rsci_idat;
  reg [15:0] out1_rsci_idat;
  reg out1_rsc_triosy_obj_ld;
  reg main_stage_0_3;
  reg reg_in1_rsc_triosy_obj_ld_cse;
  reg [15:0] regs_1_sva;
  reg [15:0] regs_0_sva;
  reg [15:0] MAC_asn_itm;
  reg [15:0] MAC_asn_62_itm;
  reg [15:0] MAC_asn_64_itm;
  reg [15:0] MAC_asn_65_itm;
  reg [15:0] MAC_asn_66_itm;
  reg [15:0] MAC_asn_67_itm;
  reg [15:0] MAC_asn_68_itm;
  reg [15:0] MAC_asn_69_itm;
  reg [15:0] MAC_asn_70_itm;
  reg [15:0] MAC_asn_71_itm;
  reg [15:0] MAC_asn_72_itm;
  reg [15:0] MAC_asn_73_itm;
  reg [15:0] MAC_asn_74_itm;
  reg [15:0] MAC_asn_75_itm;
  reg [15:0] MAC_asn_76_itm;
  reg [15:0] MAC_asn_77_itm;
  reg [15:0] MAC_asn_78_itm;
  reg [15:0] MAC_asn_79_itm;
  reg [15:0] MAC_asn_80_itm;
  reg [15:0] MAC_asn_81_itm;
  reg [15:0] MAC_asn_82_itm;
  reg [15:0] MAC_asn_83_itm;
  reg [15:0] MAC_asn_84_itm;
  reg [15:0] MAC_asn_85_itm;
  reg [15:0] MAC_asn_86_itm;
  reg [15:0] MAC_asn_87_itm;
  reg [15:0] MAC_asn_88_itm;
  reg [15:0] MAC_asn_89_itm;
  reg [15:0] MAC_asn_90_itm;
  reg [29:0] MAC_1_mul_itm_1;
  wire signed [32:0] nl_MAC_1_mul_itm_1;
  reg [29:0] MAC_2_mul_itm_1;
  wire signed [32:0] nl_MAC_2_mul_itm_1;
  reg [29:0] MAC_3_mul_itm_1;
  wire signed [32:0] nl_MAC_3_mul_itm_1;
  reg [29:0] MAC_4_mul_itm_1;
  wire signed [32:0] nl_MAC_4_mul_itm_1;
  reg [29:0] MAC_5_mul_itm_1;
  wire signed [32:0] nl_MAC_5_mul_itm_1;
  reg [29:0] MAC_6_mul_itm_1;
  wire signed [32:0] nl_MAC_6_mul_itm_1;
  reg [29:0] MAC_7_mul_itm_1;
  wire signed [32:0] nl_MAC_7_mul_itm_1;
  reg [29:0] MAC_8_mul_itm_1;
  wire signed [32:0] nl_MAC_8_mul_itm_1;
  reg [29:0] MAC_acc_17_itm_1;
  wire [30:0] nl_MAC_acc_17_itm_1;
  reg [29:0] MAC_9_mul_itm_1;
  wire signed [32:0] nl_MAC_9_mul_itm_1;
  reg [29:0] MAC_10_mul_itm_1;
  wire signed [32:0] nl_MAC_10_mul_itm_1;
  reg [29:0] MAC_11_mul_itm_1;
  wire signed [32:0] nl_MAC_11_mul_itm_1;
  reg [29:0] MAC_12_mul_itm_1;
  wire signed [32:0] nl_MAC_12_mul_itm_1;
  reg [29:0] MAC_13_mul_itm_1;
  wire signed [32:0] nl_MAC_13_mul_itm_1;
  reg [29:0] MAC_14_mul_itm_1;
  wire signed [32:0] nl_MAC_14_mul_itm_1;
  reg [29:0] MAC_15_mul_itm_1;
  wire signed [32:0] nl_MAC_15_mul_itm_1;
  reg [29:0] MAC_16_mul_itm_1;
  wire signed [32:0] nl_MAC_16_mul_itm_1;
  reg [29:0] MAC_acc_itm_1;
  wire [30:0] nl_MAC_acc_itm_1;

  wire[29:0] MAC_16_acc_2_nl;
  wire[30:0] nl_MAC_16_acc_2_nl;
  wire[29:0] MAC_acc_15_nl;
  wire[30:0] nl_MAC_acc_15_nl;
  wire[29:0] MAC_acc_11_nl;
  wire[30:0] nl_MAC_acc_11_nl;
  wire[29:0] MAC_acc_10_nl;
  wire[30:0] nl_MAC_acc_10_nl;
  wire[29:0] MAC_acc_14_nl;
  wire[30:0] nl_MAC_acc_14_nl;
  wire[29:0] MAC_acc_9_nl;
  wire[30:0] nl_MAC_acc_9_nl;
  wire[29:0] MAC_acc_8_nl;
  wire[30:0] nl_MAC_acc_8_nl;
  wire[29:0] MAC_acc_13_nl;
  wire[30:0] nl_MAC_acc_13_nl;
  wire[29:0] MAC_acc_7_nl;
  wire[30:0] nl_MAC_acc_7_nl;
  wire[29:0] MAC_acc_6_nl;
  wire[30:0] nl_MAC_acc_6_nl;
  wire[29:0] MAC_acc_16_nl;
  wire[30:0] nl_MAC_acc_16_nl;
  wire[29:0] MAC_acc_5_nl;
  wire[30:0] nl_MAC_acc_5_nl;
  wire[29:0] MAC_acc_12_nl;
  wire[30:0] nl_MAC_acc_12_nl;
  wire[16:0] MAC_9_acc_3_nl;
  wire[17:0] nl_MAC_9_acc_3_nl;
  wire[16:0] MAC_10_acc_3_nl;
  wire[17:0] nl_MAC_10_acc_3_nl;
  wire[16:0] MAC_11_acc_3_nl;
  wire[17:0] nl_MAC_11_acc_3_nl;
  wire[16:0] MAC_12_acc_3_nl;
  wire[17:0] nl_MAC_12_acc_3_nl;
  wire[16:0] MAC_13_acc_3_nl;
  wire[17:0] nl_MAC_13_acc_3_nl;
  wire[16:0] MAC_14_acc_3_nl;
  wire[17:0] nl_MAC_14_acc_3_nl;
  wire[16:0] MAC_15_acc_3_nl;
  wire[17:0] nl_MAC_15_acc_3_nl;
  wire[16:0] MAC_16_acc_3_nl;
  wire[17:0] nl_MAC_16_acc_3_nl;
  wire[16:0] MAC_1_acc_3_nl;
  wire[17:0] nl_MAC_1_acc_3_nl;
  wire[16:0] MAC_2_acc_3_nl;
  wire[17:0] nl_MAC_2_acc_3_nl;
  wire[16:0] MAC_3_acc_3_nl;
  wire[17:0] nl_MAC_3_acc_3_nl;
  wire[16:0] MAC_4_acc_3_nl;
  wire[17:0] nl_MAC_4_acc_3_nl;
  wire[16:0] MAC_5_acc_3_nl;
  wire[17:0] nl_MAC_5_acc_3_nl;
  wire[16:0] MAC_6_acc_3_nl;
  wire[17:0] nl_MAC_6_acc_3_nl;
  wire[16:0] MAC_7_acc_3_nl;
  wire[17:0] nl_MAC_7_acc_3_nl;
  wire[16:0] MAC_8_acc_3_nl;
  wire[17:0] nl_MAC_8_acc_3_nl;

  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_v2 #(.rscid(32'sd1),
  .width(32'sd512)) coeffs_rsci (
      .d(coeffs_rsci_d),
      .z(coeffs_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd16)) in1_rsci (
      .dat(in1_rsc_dat),
      .idat(in1_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd16)) out1_rsci (
      .idat(out1_rsci_idat),
      .dat(out1_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) coeffs_rsc_triosy_obj (
      .ld(reg_in1_rsc_triosy_obj_ld_cse),
      .lz(coeffs_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) in1_rsc_triosy_obj (
      .ld(reg_in1_rsc_triosy_obj_ld_cse),
      .lz(in1_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) out1_rsc_triosy_obj (
      .ld(out1_rsc_triosy_obj_ld),
      .lz(out1_rsc_triosy_lz)
    );
  always @(posedge clk) begin
    if ( rst ) begin
      out1_rsc_triosy_obj_ld <= 1'b0;
      MAC_acc_17_itm_1 <= 30'b000000000000000000000000000000;
      MAC_acc_itm_1 <= 30'b000000000000000000000000000000;
      reg_in1_rsc_triosy_obj_ld_cse <= 1'b0;
      main_stage_0_3 <= 1'b0;
      MAC_9_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_10_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_11_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_12_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_13_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_14_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_15_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_16_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_1_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_2_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_3_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_4_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_5_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_6_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_7_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_8_mul_itm_1 <= 30'b000000000000000000000000000000;
      MAC_asn_89_itm <= 16'b0000000000000000;
      MAC_asn_90_itm <= 16'b0000000000000000;
      MAC_asn_87_itm <= 16'b0000000000000000;
      MAC_asn_88_itm <= 16'b0000000000000000;
      MAC_asn_85_itm <= 16'b0000000000000000;
      MAC_asn_86_itm <= 16'b0000000000000000;
      MAC_asn_83_itm <= 16'b0000000000000000;
      MAC_asn_84_itm <= 16'b0000000000000000;
      MAC_asn_81_itm <= 16'b0000000000000000;
      MAC_asn_82_itm <= 16'b0000000000000000;
      MAC_asn_79_itm <= 16'b0000000000000000;
      MAC_asn_80_itm <= 16'b0000000000000000;
      MAC_asn_77_itm <= 16'b0000000000000000;
      MAC_asn_78_itm <= 16'b0000000000000000;
      MAC_asn_75_itm <= 16'b0000000000000000;
      MAC_asn_76_itm <= 16'b0000000000000000;
      MAC_asn_73_itm <= 16'b0000000000000000;
      MAC_asn_74_itm <= 16'b0000000000000000;
      MAC_asn_71_itm <= 16'b0000000000000000;
      MAC_asn_72_itm <= 16'b0000000000000000;
      MAC_asn_69_itm <= 16'b0000000000000000;
      MAC_asn_70_itm <= 16'b0000000000000000;
      MAC_asn_67_itm <= 16'b0000000000000000;
      MAC_asn_68_itm <= 16'b0000000000000000;
      MAC_asn_65_itm <= 16'b0000000000000000;
      MAC_asn_66_itm <= 16'b0000000000000000;
      MAC_asn_itm <= 16'b0000000000000000;
      regs_1_sva <= 16'b0000000000000000;
      MAC_asn_64_itm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
      MAC_asn_62_itm <= 16'b0000000000000000;
    end
    else begin
      out1_rsc_triosy_obj_ld <= main_stage_0_3;
      MAC_acc_17_itm_1 <= nl_MAC_acc_17_itm_1[29:0];
      MAC_acc_itm_1 <= nl_MAC_acc_itm_1[29:0];
      reg_in1_rsc_triosy_obj_ld_cse <= 1'b1;
      main_stage_0_3 <= reg_in1_rsc_triosy_obj_ld_cse;
      MAC_9_mul_itm_1 <= nl_MAC_9_mul_itm_1[29:0];
      MAC_10_mul_itm_1 <= nl_MAC_10_mul_itm_1[29:0];
      MAC_11_mul_itm_1 <= nl_MAC_11_mul_itm_1[29:0];
      MAC_12_mul_itm_1 <= nl_MAC_12_mul_itm_1[29:0];
      MAC_13_mul_itm_1 <= nl_MAC_13_mul_itm_1[29:0];
      MAC_14_mul_itm_1 <= nl_MAC_14_mul_itm_1[29:0];
      MAC_15_mul_itm_1 <= nl_MAC_15_mul_itm_1[29:0];
      MAC_16_mul_itm_1 <= nl_MAC_16_mul_itm_1[29:0];
      MAC_1_mul_itm_1 <= nl_MAC_1_mul_itm_1[29:0];
      MAC_2_mul_itm_1 <= nl_MAC_2_mul_itm_1[29:0];
      MAC_3_mul_itm_1 <= nl_MAC_3_mul_itm_1[29:0];
      MAC_4_mul_itm_1 <= nl_MAC_4_mul_itm_1[29:0];
      MAC_5_mul_itm_1 <= nl_MAC_5_mul_itm_1[29:0];
      MAC_6_mul_itm_1 <= nl_MAC_6_mul_itm_1[29:0];
      MAC_7_mul_itm_1 <= nl_MAC_7_mul_itm_1[29:0];
      MAC_8_mul_itm_1 <= nl_MAC_8_mul_itm_1[29:0];
      MAC_asn_89_itm <= MAC_asn_87_itm;
      MAC_asn_90_itm <= MAC_asn_89_itm;
      MAC_asn_87_itm <= MAC_asn_85_itm;
      MAC_asn_88_itm <= MAC_asn_90_itm;
      MAC_asn_85_itm <= MAC_asn_83_itm;
      MAC_asn_86_itm <= MAC_asn_88_itm;
      MAC_asn_83_itm <= MAC_asn_81_itm;
      MAC_asn_84_itm <= MAC_asn_86_itm;
      MAC_asn_81_itm <= MAC_asn_79_itm;
      MAC_asn_82_itm <= MAC_asn_84_itm;
      MAC_asn_79_itm <= MAC_asn_77_itm;
      MAC_asn_80_itm <= MAC_asn_82_itm;
      MAC_asn_77_itm <= MAC_asn_75_itm;
      MAC_asn_78_itm <= MAC_asn_80_itm;
      MAC_asn_75_itm <= MAC_asn_73_itm;
      MAC_asn_76_itm <= MAC_asn_78_itm;
      MAC_asn_73_itm <= MAC_asn_71_itm;
      MAC_asn_74_itm <= MAC_asn_76_itm;
      MAC_asn_71_itm <= MAC_asn_69_itm;
      MAC_asn_72_itm <= MAC_asn_74_itm;
      MAC_asn_69_itm <= MAC_asn_67_itm;
      MAC_asn_70_itm <= MAC_asn_72_itm;
      MAC_asn_67_itm <= MAC_asn_65_itm;
      MAC_asn_68_itm <= MAC_asn_70_itm;
      MAC_asn_65_itm <= regs_1_sva;
      MAC_asn_66_itm <= MAC_asn_68_itm;
      MAC_asn_itm <= MAC_asn_62_itm;
      regs_1_sva <= regs_0_sva;
      MAC_asn_64_itm <= MAC_asn_66_itm;
      regs_0_sva <= in1_rsci_idat;
      MAC_asn_62_itm <= MAC_asn_64_itm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out1_rsci_idat <= 16'b0000000000000000;
    end
    else if ( main_stage_0_3 ) begin
      out1_rsci_idat <= readslicef_30_16_14((MAC_16_acc_2_nl));
    end
  end
  assign nl_MAC_acc_11_nl = MAC_1_mul_itm_1 + MAC_2_mul_itm_1;
  assign MAC_acc_11_nl = nl_MAC_acc_11_nl[29:0];
  assign nl_MAC_acc_10_nl = MAC_3_mul_itm_1 + MAC_4_mul_itm_1;
  assign MAC_acc_10_nl = nl_MAC_acc_10_nl[29:0];
  assign nl_MAC_acc_15_nl = (MAC_acc_11_nl) + (MAC_acc_10_nl);
  assign MAC_acc_15_nl = nl_MAC_acc_15_nl[29:0];
  assign nl_MAC_acc_9_nl = MAC_5_mul_itm_1 + MAC_6_mul_itm_1;
  assign MAC_acc_9_nl = nl_MAC_acc_9_nl[29:0];
  assign nl_MAC_acc_8_nl = MAC_7_mul_itm_1 + MAC_8_mul_itm_1;
  assign MAC_acc_8_nl = nl_MAC_acc_8_nl[29:0];
  assign nl_MAC_acc_14_nl = (MAC_acc_9_nl) + (MAC_acc_8_nl);
  assign MAC_acc_14_nl = nl_MAC_acc_14_nl[29:0];
  assign nl_MAC_acc_17_itm_1  = (MAC_acc_15_nl) + (MAC_acc_14_nl);
  assign nl_MAC_acc_7_nl = MAC_9_mul_itm_1 + MAC_10_mul_itm_1;
  assign MAC_acc_7_nl = nl_MAC_acc_7_nl[29:0];
  assign nl_MAC_acc_6_nl = MAC_11_mul_itm_1 + MAC_12_mul_itm_1;
  assign MAC_acc_6_nl = nl_MAC_acc_6_nl[29:0];
  assign nl_MAC_acc_13_nl = (MAC_acc_7_nl) + (MAC_acc_6_nl);
  assign MAC_acc_13_nl = nl_MAC_acc_13_nl[29:0];
  assign nl_MAC_acc_5_nl = MAC_13_mul_itm_1 + MAC_14_mul_itm_1;
  assign MAC_acc_5_nl = nl_MAC_acc_5_nl[29:0];
  assign nl_MAC_acc_12_nl = MAC_15_mul_itm_1 + MAC_16_mul_itm_1;
  assign MAC_acc_12_nl = nl_MAC_acc_12_nl[29:0];
  assign nl_MAC_acc_16_nl = (MAC_acc_5_nl) + (MAC_acc_12_nl);
  assign MAC_acc_16_nl = nl_MAC_acc_16_nl[29:0];
  assign nl_MAC_acc_itm_1  = (MAC_acc_13_nl) + (MAC_acc_16_nl);
  assign nl_MAC_9_acc_3_nl = conv_s2s_16_17(MAC_asn_75_itm) + conv_s2s_16_17(MAC_asn_76_itm);
  assign MAC_9_acc_3_nl = nl_MAC_9_acc_3_nl[16:0];
  assign nl_MAC_9_mul_itm_1  = $signed((MAC_9_acc_3_nl)) * $signed((coeffs_rsci_d[143:128]));
  assign nl_MAC_10_acc_3_nl = conv_s2s_16_17(MAC_asn_77_itm) + conv_s2s_16_17(MAC_asn_78_itm);
  assign MAC_10_acc_3_nl = nl_MAC_10_acc_3_nl[16:0];
  assign nl_MAC_10_mul_itm_1  = $signed((MAC_10_acc_3_nl)) * $signed((coeffs_rsci_d[159:144]));
  assign nl_MAC_11_acc_3_nl = conv_s2s_16_17(MAC_asn_79_itm) + conv_s2s_16_17(MAC_asn_80_itm);
  assign MAC_11_acc_3_nl = nl_MAC_11_acc_3_nl[16:0];
  assign nl_MAC_11_mul_itm_1  = $signed((MAC_11_acc_3_nl)) * $signed((coeffs_rsci_d[175:160]));
  assign nl_MAC_12_acc_3_nl = conv_s2s_16_17(MAC_asn_81_itm) + conv_s2s_16_17(MAC_asn_82_itm);
  assign MAC_12_acc_3_nl = nl_MAC_12_acc_3_nl[16:0];
  assign nl_MAC_12_mul_itm_1  = $signed((MAC_12_acc_3_nl)) * $signed((coeffs_rsci_d[191:176]));
  assign nl_MAC_13_acc_3_nl = conv_s2s_16_17(MAC_asn_83_itm) + conv_s2s_16_17(MAC_asn_84_itm);
  assign MAC_13_acc_3_nl = nl_MAC_13_acc_3_nl[16:0];
  assign nl_MAC_13_mul_itm_1  = $signed((MAC_13_acc_3_nl)) * $signed((coeffs_rsci_d[207:192]));
  assign nl_MAC_14_acc_3_nl = conv_s2s_16_17(MAC_asn_85_itm) + conv_s2s_16_17(MAC_asn_86_itm);
  assign MAC_14_acc_3_nl = nl_MAC_14_acc_3_nl[16:0];
  assign nl_MAC_14_mul_itm_1  = $signed((MAC_14_acc_3_nl)) * $signed((coeffs_rsci_d[223:208]));
  assign nl_MAC_15_acc_3_nl = conv_s2s_16_17(MAC_asn_87_itm) + conv_s2s_16_17(MAC_asn_88_itm);
  assign MAC_15_acc_3_nl = nl_MAC_15_acc_3_nl[16:0];
  assign nl_MAC_15_mul_itm_1  = $signed((MAC_15_acc_3_nl)) * $signed((coeffs_rsci_d[239:224]));
  assign nl_MAC_16_acc_3_nl = conv_s2s_16_17(MAC_asn_89_itm) + conv_s2s_16_17(MAC_asn_90_itm);
  assign MAC_16_acc_3_nl = nl_MAC_16_acc_3_nl[16:0];
  assign nl_MAC_16_mul_itm_1  = $signed((MAC_16_acc_3_nl)) * $signed((coeffs_rsci_d[255:240]));
  assign nl_MAC_1_acc_3_nl = conv_s2s_16_17(in1_rsci_idat) + conv_s2s_16_17(MAC_asn_itm);
  assign MAC_1_acc_3_nl = nl_MAC_1_acc_3_nl[16:0];
  assign nl_MAC_1_mul_itm_1  = $signed((MAC_1_acc_3_nl)) * $signed((coeffs_rsci_d[15:0]));
  assign nl_MAC_2_acc_3_nl = conv_s2s_16_17(regs_0_sva) + conv_s2s_16_17(MAC_asn_62_itm);
  assign MAC_2_acc_3_nl = nl_MAC_2_acc_3_nl[16:0];
  assign nl_MAC_2_mul_itm_1  = $signed((MAC_2_acc_3_nl)) * $signed((coeffs_rsci_d[31:16]));
  assign nl_MAC_3_acc_3_nl = conv_s2s_16_17(regs_1_sva) + conv_s2s_16_17(MAC_asn_64_itm);
  assign MAC_3_acc_3_nl = nl_MAC_3_acc_3_nl[16:0];
  assign nl_MAC_3_mul_itm_1  = $signed((MAC_3_acc_3_nl)) * $signed((coeffs_rsci_d[47:32]));
  assign nl_MAC_4_acc_3_nl = conv_s2s_16_17(MAC_asn_65_itm) + conv_s2s_16_17(MAC_asn_66_itm);
  assign MAC_4_acc_3_nl = nl_MAC_4_acc_3_nl[16:0];
  assign nl_MAC_4_mul_itm_1  = $signed((MAC_4_acc_3_nl)) * $signed((coeffs_rsci_d[63:48]));
  assign nl_MAC_5_acc_3_nl = conv_s2s_16_17(MAC_asn_67_itm) + conv_s2s_16_17(MAC_asn_68_itm);
  assign MAC_5_acc_3_nl = nl_MAC_5_acc_3_nl[16:0];
  assign nl_MAC_5_mul_itm_1  = $signed((MAC_5_acc_3_nl)) * $signed((coeffs_rsci_d[79:64]));
  assign nl_MAC_6_acc_3_nl = conv_s2s_16_17(MAC_asn_69_itm) + conv_s2s_16_17(MAC_asn_70_itm);
  assign MAC_6_acc_3_nl = nl_MAC_6_acc_3_nl[16:0];
  assign nl_MAC_6_mul_itm_1  = $signed((MAC_6_acc_3_nl)) * $signed((coeffs_rsci_d[95:80]));
  assign nl_MAC_7_acc_3_nl = conv_s2s_16_17(MAC_asn_71_itm) + conv_s2s_16_17(MAC_asn_72_itm);
  assign MAC_7_acc_3_nl = nl_MAC_7_acc_3_nl[16:0];
  assign nl_MAC_7_mul_itm_1  = $signed((MAC_7_acc_3_nl)) * $signed((coeffs_rsci_d[111:96]));
  assign nl_MAC_8_acc_3_nl = conv_s2s_16_17(MAC_asn_73_itm) + conv_s2s_16_17(MAC_asn_74_itm);
  assign MAC_8_acc_3_nl = nl_MAC_8_acc_3_nl[16:0];
  assign nl_MAC_8_mul_itm_1  = $signed((MAC_8_acc_3_nl)) * $signed((coeffs_rsci_d[127:112]));
  assign nl_MAC_16_acc_2_nl = MAC_acc_17_itm_1 + MAC_acc_itm_1;
  assign MAC_16_acc_2_nl = nl_MAC_16_acc_2_nl[29:0];

  function automatic [15:0] readslicef_30_16_14;
    input [29:0] vector;
    reg [29:0] tmp;
  begin
    tmp = vector >> 14;
    readslicef_30_16_14 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] conv_s2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_17 = {vector[15], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, coeffs_rsc_z, coeffs_rsc_triosy_lz, in1_rsc_dat, in1_rsc_triosy_lz, out1_rsc_dat,
      out1_rsc_triosy_lz
);
  input clk;
  input rst;
  input [511:0] coeffs_rsc_z;
  output coeffs_rsc_triosy_lz;
  input [15:0] in1_rsc_dat;
  output in1_rsc_triosy_lz;
  output [15:0] out1_rsc_dat;
  output out1_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .coeffs_rsc_z(coeffs_rsc_z),
      .coeffs_rsc_triosy_lz(coeffs_rsc_triosy_lz),
      .in1_rsc_dat(in1_rsc_dat),
      .in1_rsc_triosy_lz(in1_rsc_triosy_lz),
      .out1_rsc_dat(out1_rsc_dat),
      .out1_rsc_triosy_lz(out1_rsc_triosy_lz)
    );
endmodule



